`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
n1ZuUH2dirbOUNmJGmvhFxEwWX8lUoW7BrrVEG7L0mTqB5eIuFo364LJkdRIF7EQcbR6uiIy+RiH
y0D5ieFc1Q==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Kutl0if69rIr24Z7o8dj8aUUlKMGnUUhvd2udyrnvwBpvFNHNwZl5EN9+pwQZAkI3cDBNF5pU1gw
vOkuyefEh9+JvIqwB3xdPqsZGTVjipLzn4JRo4SxzaGZlmmaLpgaS9STCvNckcFkDhkynzLi+Ehv
lk+1bhCHPsUmgdTXiCA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FmvxmF+VX/0t4G5E327myocynnZApSzZMLk4o+oh7IJVWp9j0r1BZDLvHGFzpBXuSG3pKE6UEC3r
xhRO8XeU+DpZSfeio27OAiZn+nB8IWZ+qMUzo+6CxvQddxDDpdGMdTwXiQ6eELK2s6dk5AZnezBh
rD1dapvR4d9M/dWBdD8QvkCkES2yAEUcddgaz67GOe1TiQQTwQjseKKk46qTrlJJ4s23J/hFenVP
mYxtHPL8WDA2WinOCyvALtIH01n7pT+24PQwmzN0Sc6zhsP8C06U92ESVBQS4NDeQ0jW1F76ORaE
xylXFzcIHjgGeDNq3UoVEnMjpqSiKgTvy/V1Rw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tGyaBXN77jWulBSnKXpxTSD4pLuUs2u22mUdHwaIBjLQH0xGziSLGR4W0lgB7eMVsZLeFS104Ahc
1pHoakxmGRyT0bjFRHsr0DVKvxRYKoDZLuxTxAAsVKUy3AICMhhgqsej3qtEmvBjLDSJhpu2wUiR
jM//wf3t1sp732/2mUIcWaTEMRTd/e/KrpDjno48dZf8HFtDVoxdBAUWVvodoDMc3HYjwvsvo0z3
YoFMpAIkxf5nz5c2n7JKHEndy/Wd8uTz2Zaeir2MEkj0iLBQpQ3qLIKHWd9AKU7MuaVfFunBNy/F
Fojm0cTSOxfAC/6DrAdBW1QrIHDohQod+FeREA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CxKo2EOwQBx0vCD9C+mxwnn2l8PHkpwuyQ3G1DmSUwaD6PCV6tI70ERrLREXoeUhlQiQblEH10UR
+PsxiYshLY3Nq3JPgB1qRiLKR1MjIKk1yBSt/0ka7Fx4n7U10QvEgElO7ETG2x9lr5d33Ud3LrRG
VSwxXUXfYLLsLcyH0cUm6qwYufbGl5G/N7XAPsTZvZ86kUW02UpLLuDrPLFSrymX52PEhjPXbTjx
pPs16R3CqbXtcfq2LKDYLLrVXsEzRydjilnaST0QoJiXaF8LKysVA02qKfMUDZLY8cGNMh8Pmttj
ZrVcomrVWyZYU4quuJoFY9yXgw8RubLa9Wbrnw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jWM1ZcUZ1AYMmY6i+gHD4c6V5YfJmFGSK14V7L1POJQgY3BNt6qiIrv6J38koIgetYmAJXdIwDPP
x/Jcf3eSO+bRJ/V3oDwpbYE4XTHTFA/KO3LsN/PKB6GB9jdlGBUamFkkZDvlnsPwnz2q699fi3+d
e5AShX4PFBcWkGWgZj0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jkA40ENH9mZ0YnNeJuJ65aFhaT0NJQ8OriHpHpzE+Gg1eR/0re8Au2TmtTJhDUyoP6QjY9UwCUxt
4MhGJQhVgC/pwOP84HJ8DFnxoJRQ4oe46OeepGKasVYSCtlkGFrpjV1JJd3S/m4we3snN5ab2PHK
Xc9CSeL6tnB4fwQAsveTO99yD6KD9jjW1ndrpSJJwCRJ0HNpSp5IYvIwT1iIlBtd8KyVl6lKIsr1
qw7JuUNywF1UmlYgKVqaf+tN5BCtCDkOqhl5VG3SSH0OiiC1uNkgULPYu1mPUYxHVwAWRQFQwxDQ
bpraZPSoIK2cReAv8n5pTnL1cOcSxM3hGBb7rg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 55552)
`protect data_block
4DJiChpKpziauk5p+z+vJ3k3nV+cBCcjMhUWuy4ovUJYdhqMjqYWXwUCgpbiewEIQaiojGXnlMop
A4xHNa9IryC3v0uvtheyuhZoeyvKeIYj5D15sMDvDPKe4igPUups5jX49WJvxNpWX0WUw3tamLIt
NWByfjVJAWjB6b4BOtWft1pSHfvCbl68bqYi6I9dwwJYAmW3VoP3o82GTRluvpeEGnBW3jgQCxSb
EymRV4OntUfVcl5KL8epZTMx8xUxMRuTMyomVjsj/3mzUJq2y+5OZZFzaTiDjmFn5WTKeZuVtZio
mlpNvCjvPWdDoQ+J5Y22NTicwuXpifmULwNHKl1L7IqarBAKebNLrozJdDj/TpwQX+/8YRvOcQWZ
o6bXwG5/DhlFMwYGrXa0pV1K47mKb7fzgGFh3UT+ZLNvPVrwWxy6Chei3DqA0ZZlFiIXl8pqRE2t
sp1vvMyywmKmvUBKPMOfYTPNSDYThxri1rpeWLi4qj9qR4EIx7WNhfwBtFYs1yffmgvGI/xcvQF6
EJFrDVDpQ3wfWC0SWzwFs/+0Y++O1tNHhrRQ0VrQOBwzddZVrEI5y9mOn7YR/s555Qx/2YEXh56I
RwxEBA7Y1GZpInr4n/Zq+6lBCs9gmVmoneyuV7xxAPN3FXFEawwgmiezZl8uF5MGYFjTIch+bpnZ
XCedvjRnQ4xcSqgE9zlAhVrt1WNceAOTDSoDJUqog9ZCMq0dcV7RhSTa1tmv28reHpJz9KIQS38I
T2VXU3/KHJqvPwtXmp92Gg7R2SnafnZBiF8MaX2YvojhOfO7J1gjaqp/dHMcjFMX3+Wx8OfrlUNY
juDJLhxUsV5OFp3Z3UvPpS3+5hWy0NbeUU1lA9TywDoAuartYSdAX/OLHr4tZ9/TM/9V0mzDzOOq
1B2fDLace0CzpTdFWjbJbq5/MvMbJaHWTG90o0vyhoEZ1f0x+BVkUpVJSznYVLycKjx8WHuSzqzH
09jrF97N9LlLu/qdYIlEl7K0hBTscdbUUWMAjgByKR+STn+MNklsZzjj87fFbY9ziU2+Oyn1We/m
cY6vmqFvrq+tf0DwkoriXE8+Youvb1/boAbIuMHoFrxfYj0TvSTThMzdKrbwZBQpEozzgdWDNAU2
LdvopKryrNYMauOlc5L0pkbuWukhr2urQx3EIiHgXwK6mPNBWwe1kcGQCXmGwFAvtLtc68+GLYUt
9yVpU2a5lt4IKT5jnpB1oHY4+KvY1AUc71nECIot0r9wSElkWDI4+esVYLoSABAKnuas2as7YsKb
W5pwcS4lzsQ3xWVUgHhZSRwDMRCEvAI9+WA44hag9Gev8TGYM2BTOhK8CXPqdIgR67KEZnAk/259
sqExoZDBdXOwyBxyYfUmlx0AqdQ2ZVxeucPZJ9oO/4U58+B7N7JSwFv7KE6NcuYOK3Hq/JNZbOSZ
9Rf6G0lfSxNaKOzXx24yAGAAV9Yq7OHrKeYHS3myWMl0y3VM22Q3R8DaFL5/hli+6a2Uhaygl7N2
lQB8A9StEdW9quE6b4CfemqqCb5l9PzZlAaFhPFPBtpOZYo/8N4lga39nj1iSeuhLJ/dJkarl8NM
yn9xEg9YRFObF5XmHuPPa7lHQ1yruNO+G1vXzHGrCW/YrQgal7Ot/9Suvgy3T9y98F+8q1GHQSbM
WMwKOGXR5oY2Ajd3I93i7XKJKBjv9uGia+5KAuhNhb/VXqmb/p1SdVWH1ExH3tOFG7CU31iwkwbq
JfJADVwcV8BkfJGNJugSdZAuo3CRftpEukoaYV+tNv1C34btfg+N+VZouBJ7bgpvdnsylU2rgy2u
DRl27OvcQ0WZHZtVyqMURHMQasMNYcWgfYt+ZmumVErOd496TmWvtwGfBrQM0ZSOtFOL4STyg14w
1NCyqkph81E5t3cI3C6lyY+l3rn9ziDyX5naue9VCiVByPeshddBlB1hOw1LpESoqyU14T3g8A+C
rKBsKQE8i9dHWGVXk2eUlEv6pUBBXD5BBFGSRfnmuHkngrmkGO0OzAl2zjPKuMEWMvBiHiTjDXYb
/o9vJu+MlwJZAuIgQ4tVGjrlbDHamjfg+OOWox1oMT3LsemR9MIa69yvOMlE+ESa+mfcZAb8JEid
sMKjZ8IagjA/qia4ngl8VPwdEIYkEMBrvOMNVs8ehgvNjeeTu5xlS2S3Ic3vGt3FaJlE+JcPrYEP
3jCBgJIKKl8fE/gjV4emMXt7ETrgqkKnlgnRpr7IRcxoh9OYTX3t6Kkj1yOtDNmrqJl9Eagcnwm/
7jrCqsCBy0d5U0b6ZmjZatPm5d1lN29mL/hI+Ngwiw/xztvzUtoFD56XxfNZmcxVuEfQURMqT5Xn
xLsxE/O9kj+g4mH/GNnpgziOJr0Uww0dxiTvzcGng2+88zkcFwhkkqKwSzPkJQuV2HMW4bwghzWz
oHFqz1CT15TpH0xkw/7hsqIonjnpln0O4YfPbAg42mqcTeJ1T7UCsdTchanUUzPiKrtFZWnhs4jD
HY7Us2igT4K85fGQ2TXhmlhlcREyd4iy+pmH7xPh1VVNwWuyhF63JUOdcfl6oqCoiWndq26Wy03e
4uDbxJCuPes/JJjImge8SHcVWWufuAN2vJKLBJ90dy6dxH35f1gcpL8b71MdmRlWT9qBPgWpkyUK
xOf2jlXykU5/kriGlvkKE0UWB3Oof+00p2DRhp3Gwt/SeOuNpCZ3w83V3xWB3G8VFVIpoBYzBWLU
siPjVjRSUcqo97x70De0m/S4DumqR8scVdkLcr4hncQaTtXUe0E/+zyiyk6SNR5MF5BQ8bcw+XQp
4TZ8oj3wtgi5sWjzdDF569fKXkAUrtNrWF/oZfrMgL4XeC0LdrqA0rWSGuHQFum9llO2ZZCCahpM
bAP+1sz3JfXbSA6r78F8a7TCDM2GwY7twGPiV963oFPus4ZA8bk3OOPHn2OZIK4hmHTmI3FBD/Dc
cvwEbRaRIpSajK5+Qil9nFY8lM7PdVO3sZ+p2JDzf3gAJA2hR5CfHIAoko9oXq5yGpiO1EFNg/3Q
7LBJ0bjbGpFXYXcNkjnQCtfwlf4JffkW52bNCJgfe2p9omufJTir9KpYsh6wVq36a/1yh5/b1Syl
uctIc9jsel8M4N/eDZnzHi2vOO9qalf3FYMSR1h9sfuWFNz8F5LL/LDQwWLMnOSkoctHKR4Zf3ne
05+RcHtE9W65SlP5iX1kSpwsJOgSX1a3QTaA1U1kBiMaynzTdvB7NtZF6Zy4u0jzJZXePg3CANnR
yKlJ746hH3OxkFlprVh+Oo3rT6BS5zirhx0xCamAXJvdqw+ITPrn4KQvqvs3xuB/JtaMcUMB9sDi
CpJRWtSj2rF3S1+soogB9A0Bl4N+KX75UdR/rxonm10P9SiHU5hhnEUCoMyb/s1wr5fsXmqXaiVx
ObWbzlN7F58NzmbanQpmC2BGGeAwkFe9IruQDV5DiiwqGueRnItoWW3qSzWF5yZSNdqTsPSrQD8M
hhxjDIdi5a+tyY5XHu1TxFcPCXXsFiqTleGwuhQk/gQN3UTAeg/2li3y7jJck+FGNiP7IVcVjFSI
pKhcJfSfrFKzLW4aTwdQz0YoroK6oNt646XTLHsCPuGIXTgwTuLI+dpv2Xe6odw9g35fNw4wvC+5
2FrFvAKUigEJ9vrYAjWyZNkUlGETFoF4rpVumW+0074wCZ9q607UdGOXZpAPh6AY5D/fuKu6NAHc
i8cdufJs5/jVbzPncACsDbPp9VyYGHQa6xhXmI9eEMm4+9WFfOr/8OpsrumOUMBaPj04NEXbSyNG
0pC64KXkqdyEuT55OuCf0CfKjT3mTB5v0X9eMAqT3ACCqwvXZjsuKq5j+q9PBIhq/5x+iH9yI+aO
mN5rjyI/cpFc9kSc76JrGRq5Zp+1aTPwhD8V5sbfft7LgG5i9NE2veo/Cdnq+bRMaWEg1xvgc8ow
BvOyrNC6HCBzyffcb7SAGBJHLV6nVIRZg8mG2J37KsAiSaY8tDY9T+RkRjTLpbzmxqpV++TH/Ae8
HLE35zLmVi/dklAAiMYTc9ND4m+b2WDvwnj/NMrScOdjiLSgPvSDP7RD+OFNbRLWKBv4mc558ga8
YkhLJQ8s79QHEQY2Kqpau4iOQRYx6bBr2GrHL2e1ZBH2y9+GdlMNwFMjM49udlxi6LO7hW/n4mXA
uQ/h9kaWLFwNjeFANmGzhZFrzgu0+l9kfhx4H9GUpPNrbd6g4IlBdQHHkuLHRvh4KfnwTnLytTv+
vIGIECNA1+tkG59Kl0+dUFCTLqyr94Djf5jrW4BRPs9FQV7HxvaFXPO8YFJh5cMY+39d0zmuhlFT
nChRXMpCnHVkMhXFuH5anJ1/2GgWxZQe0R8YtSuctBNHjdqS9kmZY02E7DpsJVt6bzEhxk6OAvsf
RAuzegNrocHuziqiE6srTqCPXNMJeHIO8H3XMAiHVeHhnBc0teobcC2dwdMxRdZYmmvQ8yNvTsgE
o1jiCRRsyodKzH80bf8juQsEsH7kHtx3n6Aa7vcLj55+8/YeCoqc483pNhOx+U9xk0zLSmrP5bQv
GcdLc7QR2EZ0cV5JD51cbFYuxm01rahks61F77jk2UDPjh0VSlDOrX32/Q85s5k0t4wvHAuTyeBE
t/nzhjPlrhyhCRYrmLgIOEca7B76hOqi65LtYDvCIQ8FN3mci2SsBETwhmCRMaQ8kkGLBUz1g3OA
uQ4bVLesYljyVNzdg3uJVNzSwRDHSpEU9nL5uwzBWB1pgOocalvHdTOF7nW88H4Mq6Ne8YG+vXs1
QWwm6Jd9YPZWYH+gYwg/2EaQmtkSKvUEjxw4uu8nUiLxJtEXgEDrhyn1h+92d2UTPAN/24KtblBD
jbi4ta2MmS2qfirOTLrZlu5PaqRpG6QJqPSZqgSPc+dhojTJeV49lBDsjIApbbfPkc9uYA/ZcmtC
4xmeap8T+XQwweMKx+U2Dg8RKLB72X5afWbdP3lTGukfV8x9JFkQtPpeS+Ufju33hStGk1rqaW2M
Y4KCdY/iMcMYKYmSkDM1wUPlOA9z5N+swNgwWlr+Y7aUkAznBhaTOpG59NODiVJcT3LKXQZU2Re9
kMqkWM/xJjuIhepRGC/9K16YLzh137IXr/KnhHgQFZ4HSxutx9JpvbFWUyBC85U1RzGZoC8F2+r4
J8R0HxPOFAqPtgj3WFfP2FA419hiQ8vCQfGWzVo3LXVPVLvHO/Ggvem0Lshoqzbew2Qggi2jOnNJ
7UG8pNu5IqJGcNG/elWsbubkwV10V4Nfag7hcXAaq2U2JKuawKlYC1Z6cbOPq4yaMHEeovKVqBR8
knHzb37Nd8spjQgbDmU+79R7Z1mCuIq5tY1Z3vmcP5mBOMGiTcWXTe9hTrrU7nbd9pTl4loSgB0z
GGR+mC3+DGuf/SaXEb0+XBOOoUpic/BO6T3IDOltjYbh6LdRZ7VnZV0fpN59/VXMmedQPTss+wQc
9vAOJTGPHZ+vxUwlI6YE929UdR7PK/sHn1e8uBTp+Kupm90CzIs47ECsChxoCLwUkndnm0B9otIH
q52wEpezQtJOoE2z7YjFUFgerZNmnj+Xv6uPNMcaNU8DrLhVqZOZLnc9x+eHJ+3Hinqtu3OrXvnO
fPPWi4PHB7aa8DGU37Kl3f18X8DVWal0qKe377ul52CjPrQJlwGSbh6fe1Z5mpsRjQ8r6DSk/wOi
WAx6MklR3U9bVc+YXdjumH23IhVXpEyGwZmJhT9P8TWSKSnm7foGqPIXbTIOJ2Xq7T5KrXlrL7Sh
PJbWBepulisIKuoAmPow/9iZiGyIo6LcSlVnk2SBYaW/du5SroRdKTfBvLTsm0hPrDeYNslXIveP
RWRLGUgthaMEABllZD1pPWAgQOz3SfaiVetcyJ527BhtWeUn32rPUqxleXH5jP72pyn404Gk2pSK
w0Rs7zMfS3y/Gdk+b8pgsVKUKzfQLd9uPaip/s/wI+6x+Ixhmc/KhUTfLIdCNWMX13+y3v25YgoL
2XFq2l+iPsdrjxN4Rhz30kXxp7lGwa3YziUC7g0gNhMKgjaG2kRXbEVrVozcgEY0fPWZbIav2bFw
B2qI+ZI6ZwdaQF1cYKzms8sUJxrlMzHY7YjSxrfZTqY+wKsn/VscEMdV4LDDRuBeNGVnbKPFamDH
I4hm7AUZFpVVxiou8OgqSIX7i8+9gTcwLezA7uX2UagXrRlqrouKHaEvw2ATBsKUN70HncJ2jhaI
PoUbi4ayjgtkHnf1LbRS0bxklROl8YltyCwMCGQH97HjzYKX+EtPzBX4M9pIuM6MDMTd6+kYfAVy
P5g07vKBgrexAe5zg5iYOCTZP9xgA2Qf1bGIyJEA/5Sy0bDuIHBdwuqLB4cGPPNuBQ6au60RrYxC
7T2sv8g5IezXnGDEQXeQg6uU0nrSA1sMJDOd/pt5IE6E1r8Ve2j/pztKcBVb58fNsckm5tThRXoM
M2H4/gaPzQsglAIH5rFV+QZ7YkVDObJP/QZj6cT2DtUAlD7+2KXvMU66jssLH2SlXVEabuStsH92
C1kU7P0znmz9yclwj4bSfLntApJprgqYazqf03BoGkxf7vJ8euRYRzncH0mzxxSV6iVGUqZ1VgsX
HtqtlKoSjYBpS23ycQck4/dHa3pU8t9GyYM/2vAwRp8WL6BXCLFhjljW5SaiqJgF5xz4ZTDgN/G5
Nkz6THjGyydEff5Js4uIVWMHX13urQkmK5//zAKSv/As9sQOfCUsoB1g1zWrdKEOBc6hC2Z1eOmH
YNjoUfDX3/6BQHX6VI4ZFY3+UjHrwWkB7MjJtMWOPXt/fic1v4WXH005W9KnU7U4AaIl7EZSb+nJ
BBsXfQojsDeEhGbYJJW2VDfY2vhpGGOqCSTjFEShZNHzAQdS+VQeLrgZ09VQ6NG6BqHK9Rs9s8ct
GOWEKQjtOqevk+frh51eXcH/7HZfYzxqaZjiL3BD5//32yMtF/bejrEO/Bm2XH2siwmZ+Rwmm2nY
qEx5yyXCBeUdpEVoYaUeqRZwaO6yM5ueDp8QZBWjFdRH5uBVrvfblR4gB/jZXjpEO3uY/CR8Esk1
/ylioHQq2m1ylgRLA/uBqPzp4KMIEH3nRfMDP/2kxGR44nGKrVaBJ3EnyUdLNGjwB2bS551eHyeI
ZqJFxvf6NJ11XiuIeKWwHKBW/EAwlMVSciXSVuCedskiN941/8nVlL8XNe4HY3Towclg3RPWYeEY
0NDQgo7g6IziEtNzj/60TdoQy7NnFYVNSfo4Rg/duntZEsyvnij3VK3MumgK4Eq4763daB13Xh93
tC6LWZmJ+ZmeyhJtsjbpr2nSGe8No1pZbXZq3qYtpOb2N+xSMiNCC9GmhPjSrBb2ONWgyVtv46fe
tBhqqh9mLysM3GvhPqSxXJvRMK06H4tIG7YTC4Wn8XyiiYwLafMV6OmnY3ouX5gtTXvtFxDVre1o
s1a1jqN+/YKkQVd6ahyhe6piqhqddjZLH/vuUMKMkfGj5HnnqJotAwtZfdKEhTLuqE5cDKnpLdon
kjSBxmyaUGg7rdngqG+Qdxan0x5E9qEy9dxkwEiOqRvt+Mz78kk75GG66JKiOBRkmDRh3apycgBb
2hDn2i0jUpSd3XJ85ABCw8AIuSXSMjk9Fsv+zlDliOQfk5xgHQCm9UtoRFipsgDF+CVBRFrnBZXF
v3hTp9937S4VmZEBR5IuZEh6rBEj7neMyqSrwZJ32XHVlTfNucf63J/uHKIrA6IDPvu510t1lK2s
gl+ttU2AOROBVaS4E3fvxKsoKP7BQIVWhBtSkPlvMck4G0bpCDNcEmPc+dRa2EjUlc4sddm5rxb0
AUnMX53KAPRqQZ+04pxklOQ+H7UQXs93v5wOoVjaM0ej2BgUHqutzfU88bGz5ZspBWfdngWlt9KJ
gb2RblW++vNw80otgf9qid51yagTKsXCnhHSegrtt86eMt0Dkc88CCcon9ImUQ9LJEWGaqVXrwDB
thbrgOJWPvV0I+ZzzuEwMvlamerjnSvkN9r0RbwurhtJFVfFx80g1CqqwlXQwTRPYDRWPs4zm4Sg
p83eVsGTe11b6VHzW4oT/kbJpo7qkWECJQMDnFM2WqUPM6/VV9gvYDUSWBuMzcXjy3dd35RE04th
sepD+mh1WzTfo6MKUAwxkD1YT1J5sAALhPQxrP98o+sdUc/lv+V7l60irKU7hQxFIIC0/HHk3O51
vCPTSA/uJSuEaHq2KzQKzR90RiaXm9sWOhKjqOVDFH18yK6Rq4Y6cV9dgGrred7tgK/MHms7kvU1
uQt8Emg7DfMeEp9K4UFMUXKN4mHDwaUgcEpdxcJw1Cpnov/Hc143ryP5HdkGzVW/zjpOZ/1oVPh4
rnAnsE+P5chijfXb/aoWVmkp+UOXaPjJX2zRpBxaYGZUiIYqEEdVs8Fx360ImLTH3SRgPG7FPx67
QGT6bcOJiulLBtBstVwdnTxorN0eJwSURM4kMDOptpPWHFk8QZ+RIDwo1riLBuJn2VeeTpqvM/bc
bn/U9Zg6QHK+h36Z2DIMhQjiCAFeZ9QA1YOR+xqoL1MSMXMw767L1NRwjoIp7edpj2M8KDtr0BBb
X4Xe2V4I+PzIMDDnJqhhjjGmEQTHyOAR3jYesoQBZJRhjSjBGUJ/V8dZw5ErrHXsavgVxb0FfipP
HQx77dKleg9Ru/YraiA2F2MqkybDizSe1sKFBkxcB9HxkQqipOaPekAkS0QhP+rgpnjzkx3yiTMN
6fkY/kJf7c49liORycVy9rL4h+hENjBmb/JbuOgJMlRxhEJUp9lpG7DJ0N8SSPiC9sd/gDGH4tHc
JKNqVhsW+RK2q+43GMz/vSkFhmTS/Iiw0NHbRkduUmNvcpGqLSuhWQvNBH6ZTCTYlovnnQ+OGjr0
sMU/iDmJBJxKS0zcYEaQygESzqd9siRZOeCON8B1JMehoCC6rrtVpiQDNtdVkAwMvaI3embBxnU1
E4oI/FP7OumY7EJ8VFJfdnPD274+B6A/7WjPezEkOzETBkmvVH044MB3x5isQ7j0GfUcWNEgryQ5
4d4TPYg49nkI3m+HtmqQy2nlxetHSNbFxRGAwhvhQPiNk0l983WKMw6kaH7/kbtGXAwOTDhfGV5L
lViGjmLXEggC7KVSbpoHRo6k0YSuManxng4jIqDTJb8FfqpX7OR5vbTMNOlh4NIjhX5wOENtr9dh
zxqJNnuDlScJZgDwMLSfvZDENh7eVVnLuZzCfLtyLD2EIn2UeNJ9Bqns3+5ypZxO32c3MdZjMfKX
SdOt9/GHcd7IL0WLUNa8LTWTByilnOONRDrygk5Ofs2J29W4rURmgtjmrHgJXoELLPFtCuex6oUv
E489yo10te3Wjxm716ko7/HSPKBclJbujvAaNNCO8aWHAUy+7sxrh62/iRp4X+UQWoCh/3qqqtsp
Z73FVVtwypsZkd4HKCyQhtvQOKhMY67sXlQtFnFKKX4idHtrM+SuwPaNJ5YRyaMaluCGLvK6ln1P
RDDiSdH/dvK35a5xM4F61Wq9y7TVoqyZ/JNnWGc0cKv/CnEUqaQQ88wZz9EzRg6QLfdYD6foy5Ds
txRZP+Yg+I7PFkU0LswoA2ekGJyPDIPe6wG39JFuvNsIoDOrMDrlNSwvbRssp0v/nxFMRb9jiCxS
Pb2ljgKtgHLYwj/uvVGHROVF22Ew5LpVOZ92bI3hqa1Z4FBU4tnqoud4+PYI1XN3Oj9bAjX+f2SM
BiYWk4qAIf5AUdnfRdcPLUV72yS/K6CDB/4x42tIsNwsFgQ4eOGQ5+w5sX3qy7ik9G/CDq7+eLVw
W4o/TijlVUP2CMvAyul37P7813bRTQwhgoe2pDk/tb9qDwS5CLlQ3ocA5p9bMxsSrf7J0zQ3ZZH6
acjs0MVVxngd59J0a1B1qrgJ9qiW4Ef0oUBYbH4vMpRSjlHXSiP0ne8w0XC1SpPWoSwNTcupSu94
gdcN6QPAtM9Us6WzUXUhtZ6PYltc793MbPqfjGfx7HO5Epk3Kw7KgGr/bl37EG9c/FxpjUgmr5V1
Zt+YtqzAV9RuPA+XpALHyopBioTg5+00HU7cFlrdRlLSpcxCy6RkYY/5X9cf/l46Es1UNsDMz27U
lWs2mz0ngKemNL8uO5+nzFanr/fyqHqwyQzfrwbQf3+IS0RjZAXicp41qy2k52MqARtWWgQ/NrR0
EToVP1vu/oIJ430RU5Zk2LTa8A8gHALaT64k+5JQ2h3KvnmLao9foyPVh14pO2TH9TY9Z00DNxzw
/zLnvNzvKGpTh4pHk8HbDZmx0s0qsc2Bc0DeS1MSGSUXI0F93YDPuJhYatWBIGJ4iZ66fP2SJ8en
K6FzSSbBqiN65BRmekrwOgV/9ASieoQiRcdZYfUtLl+++bg1wL1gP0qvxdOUWvLJ34/AneTXfoD1
rgaNVFpndk9pmtoTKMhKnhWY6MQneuDVYqz+C/HWuDtc1Q8+WbXuR0L3WDqaCAIUjkLQZGXs7mw3
yJcCDEm0CwaY8ilm8RFZ8/jtETkWZFMRxpw/adA07oHkEQM+yODopG3TcZjcID3yRuLeTX3JngtW
91jhJCjxx4f7zW/0cujCdccKzC9cdJe7QNulmfXoZ1kF05N2iZl3klreKwN7B4byruFJS1DXbFYO
3B/6JpzzLiUf6/FwYNXlmJIYd8E1uXeFzgo8/wJeJGMXxco+Zkpi+xUkuUEwMMsoYa4c7EdX/e5V
wKouWrj1jCUDopGSNEqj5W4k8T9752vsfg1hKdxBl0aYqmsZ3O1PK9WanS1YyufcodWwFZRykzNo
M0+2z1h94yPdCfRjWebOdJWHd884udu2MVmYgfUCpausp8W8ds+5KChm48sf3elPnkWb0uXvPkhN
2IlTS9rwsioagFhTwMNA71Qm/flLR+wLO2RNn/ZTIqLLfdP1JLhsgLYvjRV6+O+MpIHqTnDlOJ7Z
xIlo7EPYDcyJ49E/aGhq3cZaF0SYrRNqKZypUxk1YLuRGM8ZPvCRT0rwxOqBdY9zjzoiaR+3w1/6
KgqlDRaNDkML8ubWttRJBsdhRUPzhdjM67jsgdnC89yFr6Czz+v8fLsv54oqD8tkv5AbxUydP+rE
bl8LKG7N8n1Unp71Sauab17+N/9kpdmfnGJMICAXMSoRGC+8EgoJEfhHx5/i0v4hb5NAHM7AlS6a
xqrV7nxrT/PJASLwZAW08xatyGBMRZzQYhc+G81FyW/cmu9iPrcpSqG7oNLESXwbLjgjf2ys/AeK
OGRCT8Kni2kNuwZSVqr/CWcoT/FbzpCij9gf5cJ2s6tfpQjPF+p/u6cDenx++TDyGHGSy2KH/c/Q
ACm3Ec7kpjrQNjP31UkgI8+TqsPcPvC38tRVAabfFnabURYlWVmM1Inw3i2aL+5+1i8++W+GrCTh
30P7beXjiX32sPa4UMqVSWcINBDfcM1r8gS7rhyb3S94IN0/87hHZf73GGKCZrnmgOtF5x0MJPe2
ARVowmgEQ0gpCB6WxXBcKMpLSD9Y4kUFA3VEK2rWBQOoymue994aIP0BZnAQjIyPDbwBDYBHXC+k
mqp5HfLgBhaqv02JjL/BOhx9yJ3PcuSVI/LK/7j5pxRFPv3D2AqwyGnqzysXURL+EZ7cHjeNp+0/
6jd24hvAylZYxpcM9KTgG3VJTwQ3+gtqZTda9JbTpFtD8ht7bycQdZ50m+Pn+DSQrF5PzOJiQfRz
QOeYxRRkZ0hEg/hSnH8dR2HGS+CbHQhn3xfycVBsKY4VtAnJ0dz3DLxdrbauzzNEat5zlhrozrQy
3cRAEtyVU0uh2qxn/ZtaW6W/kvqQJKwHzIacwjsH8Ut9THYzTFliIEJeWIN7w1hu3gZNyXR9g/yR
XOSbTZ7Q28JynXh4+792Wkp73d2XUGbYmkJ+wRtltit23tr60o4WpQYI8dIRvmKA+It4M4elEUd+
ED5YvsMaScK9iIcXnoU8fqrnTXnf6LLE0uCb93HkbAA1EMcOx6aa2OYM6H1U0VR8MBJy0FWqoIDF
119MbwdNKGWoE282qNXWosKhI+Sq8pjqS9iVnjF9y1l8bST8GQC4PFh8Iy0UkzX+liqhmW5oZxW5
Q6vHHV1NNJf1YS4kXsMtGlWrkUsMZeWBNshZwHnQK/gB8Qq9zxe1bJ8HHPeT04DVUsxxs4mKIpXv
veikLEDlu312eR9GNPy72NtNOGqEOIQU9FhGODqPXgkylRF6s9+ZSpO0dezRpWpzjGFN1jd81R89
DQeVttpcUxpBVgI7pe3D+rPYHDAwAP0+YtXZ3OT/K/lS9vOZU5C37f2yaop+PTj/cPZFoAUGjrcG
fBvjnvFi1wJ1VdkZrqODNregroQ1lyHLjZBZTLDhKVY+bj+2MGtKjUb1KwzgneDdfvnC/e2ybUWc
bGdjDOQ8/SL37qmOLvQcjoPyTWEN8nxlLRG6Ab6fgcSp8FHawg9F+paFZMGFg+6u1f6AkmuJ8oHE
3LByR/J+w+wEux/DWcDQd+Y76OGdMUOspZbOFd5ajl9Hlw6P0bGhlvNWa1zPfd8gkcPMErA9XHMq
ihjdaeTXEtmqE+Xrp3q7XEVxZ0flHBScyEj/TDP/dss+G9Qr7ZuSfTLJHqmT9SONsLSNLS9u+ZPB
MxaO1qiFlWW01a7RZAiJZ3qUrBYKC1d5y1PDWls0LGByfahgyZhAmI/sWgI/kGIIsWKWfnmvfUHn
SKcSmW5Hi96J/ScObf8vuV2rkCbyL07FXjLutdvoAaC1YOenvcI1pVO84PQlIygIV1tD1QEAjjoG
Tu/qdo1cQnkGy7zXeAVHBfhsT2h69GSIlxBlNDq+nynDimgOnRm5NbTAcY+gxITbs2726Hci7g9P
R5l8LbPJIWJ4jovjmf5jfz5C3wKE2n0xZnvnKDnjhgw2W50DMNySgIsx9NE9n/XBnopPg0nuDRvk
lvftycSsREeO+l76hyPBlbWNQ5EwaId9RWcLCvYjidA/CGGhVO6Y/QGybUAtiJ1nKO9CZ3DR3Vfd
f7cJOHTyr+kg8b5MDCrluRXsrCU6IiXmLBQXkH/iBnWKRTZ21s9LTGpqwMiz4BEHAAkWLB+Ts0Uv
/PQhEIyceJxsr3u1FyrxhL0ig5QSOReCQAhwIsRsHykdBW5+1Bx8LoXodZHHelg8hmd2HlD9Hiph
AdRkJJUPGBPdC01g7MQOkwKrwU0jsZUnfO9DEJsPa+/wMOXm2EsGsugLIYpEyZfrWbH47SjQ5jOU
l66W9ByNW4nxgM7d4pkWmmi2sxY57DROzqFPoLzHOcmT2MKOmVYInJ4m9HBuf+J6hQoLDOkwNbwQ
vKlRwLDg5RwpP/o7r95NdW0VhMcBir3fu9U5uqyOzVJDc+A4ToBbwslHO/1SXCAKtDwfA1yqWypR
k5ZFP6yTVf8YjEE36uRIiluZ/202uFPq9hfLtsOpgEm0wJNcoBJ7dgrP2RrgCywui+NAUqBWAZX7
+qL5quiQrljZK6SIWtzeRZAniVFrebdFVyYj5QaMIyiYPLYU67s3zEbe4qy4JiICiytaqhJeDrSE
aEO88TNMY/V21rjUfO/wjH8zSKZvXxUfILQwlUNcAZFH8WTsAr7pwgZvZdbDzIuP5gJ72e02dxAj
RSq1ER/LqdYUFSYf9IBEjC3a3QyP5nas+vV4wIvEKFUulPH+HVnQzXkKFuD9sQcaNok2Q1Oie5pq
vqZAfDPcYhWXrugpdRErmugSrb93qc8SB5jFW+5AkdoMOnYQYP4wSO5QVghzzzkOO7XBkacPG7tZ
vxQGMwALpd8nb87yVB3nsONw0i8ieoMPfgJQPIZ7t8g7ULz1NFLtKaUST7eyDtjiUsIWbmgtnZpq
qle4GO23RRIhPNlzUphuGE8v088K0Xbzcu+MnfiC4jlx9Ncq7xwWbTXeAwr9q8hbZz3LrtmoW32V
qvyxlM0JgYhtdeyEf9jn5vrfzLvvgjBl0ZvOAvK8pzOh1//L1MAtrTQ5nMteH+3koyGKrtUBusRv
GYrZk6aDKtDxlaJRpF47BZsyENXzCJ09SGPZKy7lgMpBayELdddirpEmkhYrZgJZnSRAbRIUt989
lLvUGyICAmzxLotLAgdMRcSYXOZ7HFZsw+X+MhNdj/IdQ7Y3VqFhM++modR5PJ26Gp9NqG8wf7WQ
TYCtlQih+ExDGujr/2tuPsX/e3hVWW8BxeQgVm2wPyknGCPAasqw6E1/731a7yWzs1YYgp5DwUYz
TeBRs5kHCs+fSWIyUhehkEb4Z72r4lwE5bqTz94yCnFWlCuKOe0nudHdCiqMqWkfI7C59Vq06oRn
m4oUx8LF7Z9Z1I7bEjX/DcH4rZxNqBtNB+526T3la7qOXrChfeBAOdBPLMK2BIyRtWcVKYBARKMP
WNCIu1V0NPsYcR/Ul8hTxPgkHIa7kqlzY9b0CbKagYN2vb6Mlr8NHYt7V0cPqKClPDngiKrzZ0lL
RuBn/65MBAN6oNZH604F8DCvZzmscUBekbYySUYiyLafLc8Cfcvc57eoHeO+YxG+uCFkXOopJw2L
XiAI/2u1PcphIbKuXVnftpP3TN/zPtKvMTIZ35uynoaF0tZ2HCSStIBduXJCVsU2KJ5qXbdRYzoT
W/1BtGNfb6GP+KoaRV+twYOtKZ1w+xdDL46gZHa2Dhh/124blbG+5081kWRJkA770DM5Ttbdymni
gXM5a6trTkM3RsW/qANt814m/YlguMrb8W2XjO/IvqW5DdSacoX0biEEUaOISLVNDfTerZezO2at
c66iFuohgin4KO8MUIlBulw9zL2YOcPxlRZX15BIWiwlm+J9iGzXN3dWPTVBfXkfbjYNFF1J+FGM
TyBNPySsWIrE6Iaih/uLlXQwocq741gtypBSqY3+hhOxYz/rG7nIPgYh3pm5gux1prLoxrJset3T
3yKxMPJYH841C5uKaj/CB3q9TlBBosXe7bGUSI3zsw9pG3rwci726Cc16jH0rASHG0U6GtQ1Fc1y
lPwA7v+xGEHBq9rLZP1IF8d8jYHC/W/7Gg/bXTNL3vANWOpidgHhi9VaDsJjdIXxELMwgDWv2T11
raeResQoeIIec+TRNkBaadrfHRCh7bDXTTTxiasbco6flzqInrGflbRAwEd6zTm3Os6FrVCZ5vqb
8MDedy8kYOKGj94Bh7RGhbvv6eQtDEV/4rk975DDetynm+naVV/x+RAZr4zhzt/PmvvqGfV2Jyf1
FeBr17i8380CGSxLmSvwiE9NEEFoNrYRXmDG640e4UwZDtWtofvTIfsGz9bgD1XastCPPKnOw7CX
3ehGpZ0KtwfSF3TKlcPf1gZhVjGqGegqPsuinboBhf3sx0Wqm6CvrJNHShiZGMLrJxHs98Zh4/ic
aPEtOwCTClvSUcr1MUo9cRMfNzKaE65uJoZ9cArXzGmlCd1F0RySmjlKektBA/UFPX68UCXydvoH
2P2CucfWhUPX3NvZtNDJ67nGet87txJo0qJvhVX8UJzLNzCi4taP+eEXGGulILhlTU8WHlrTILlf
2y4GhE79gQHbXT6ul2/ic8L9dZx0cMJ4VjcOfN4gmjuA7qcpH8jWhY8gROBupXdNWLoMv1yTJqYu
RcUXHydBhAVeLJrOGX+MQ39g6yBLO0KZ8Ezz+qo8uS2GYuLWzJ9LvDg0vbFWYXLCvF/PJ2dT1Lx/
302Y4JuAvpjsCI3PFW/tSWY6jMH9LnWOhLyTgHvyuwJ4PfBv6MHBMgR/qhcsIlOUwnT+MWjB/ZHO
gvVh9pPSgCjpeYIbT7ium2zNOYuWox9ArGqWwtpInFn1HWmCqA+8DEQNnyoyAgz8h4n2XGUJYI0V
mNlLsGCsY3ch8XxdUKFesMP9SKQU6gHlJw41cvV0k7IyTuBrk+BDSz/oz9W1JdNpDebZYzfPMfQm
ryE7r49e5trK7A2zONCkwfGAbmzMH3eq6hTNICouGBhF5ZilBfHfbsNNu/lg+Lc1KZe3Yjd6s3Pw
gCxem/BvbYxcdEHHPrvihGl840aSB5GCNYZNPp6/uKIoskAvajU2jcPWRnD0vkjF9PwzJe/qpmfh
75Fj+zprlyeWGS/kKfciDyRCPLS85DhD+XRsdPw/o1+FuMGqZncSwUhOir5MZJ9Y/X+sBspZs7hP
dYNSQ1Sp1NBIKWmySfY3Q7QTsiGm8rZUauofXzh6mDhnXTJM9x2t3ExVVf6L9OfkyYdwTsMjnapP
b/zltdVQXnMva4YkyNrArx83QkG6n+E3qac2KhcDfGTVjdwf5eEFS6WHpT/Ky9RcqwDu/cnzXjZ7
QHAHCIkcF/6ip0bRZsxcH/BFzUTuJ3/fz+yaiSYs5xxd2rtRw5WayzXuWW+EqD/DQ0zWmQAOXCN3
cneQnoP8FvXoR73kfySj8i943l++V8SROyF/LGp6k98zCB1WY10Sjxpsw1XFHh2w5sl38lCLgzhr
zJyam1q+bPjTE0TqBVYX9wDqeOFjsOA2/hvj4nXaa09mtxC/Bm/g5OtYFXDGv+KBhLW9qSXdr/ye
XOvHn/IMFzHddnyJlv4kvoBjrV8lyiPXTsU81hCsIxoaIZyz4Pwclt6RunfTiKCWOZu6QHgqI3Oz
K2CSDhjAFT5qBWqD5txlDSnlR/+0n0UOw2/UOusHqxvn/1vEYlB3CdpmUVtFEGZusEacRCxh1jF6
uitKbMPmPl7c8fO3MzKLgGisyQIjTdig7e2ZlhGfDUwAaiUPRanFKj9O31Y6j19PYoLR5GThdvXK
q+8s6vDYf9w9KdFk4hmhJ/sCLzRBgoHw+Dt4dSzbVA9kl5tdKf7MOqh3SmACaoEdwQgnX975VUs+
X1zTf2SrssIo5DTif+uLCLOltHSZe/UcX+HKAhSA3z/0BnOgeD+wC1EiJlARXLoANjmMFrGYKVtt
4zsQm3Qq8glo5qBfXfTZnvYV98Egqkpk1FyjWsiXqRUq/9EElGFZBhkFmDRHGWiqYH73xzcrXL/W
QLXr84Trh/7rvejChafrmg2bBKImkPvMgoYnIJdwxdN28pakXyaT+xlfEGm4q70J1Dx+wDV4VI/d
NhwliG1EQ9rMbFA1Cuheec4tDe2tldYlHw9saLfRZlcgDXNt7n+7W+nUB2l6ZSQNSVj7JRUZ+Z/L
+kINYNQcAKvmsi+DKuNYrswosq/JqzZFZXQNl/bRb3DYrNaC5+XvUQK8O+7hwqLF6V6wAIghnx6c
glYxURGuYu84c1l5I/VobVo1dbgd7Pb0B62lTExWpjLzK7wVasSIAool0o++ne/ePeDfPZx8RM19
L+NJv2i7q2XOXZWPpeBidTgyLGfsqFdN36spUgd+qZq7U6xMtW6+jWT4lHN8NgF+oxdLKbOTJunl
b9XFFEiLqweEqRXv8XzYPfOxgqOeHKBy495VGFcN0Z9OQ/JCRjki8VG7WUXZAijTQm4m5xWs2zBh
247X15FmbmaqdIy4OdwPtT3n0XKZr5sw2MazbRxg02NCMGAmduXr4T6cZWuz2S0a5ruDyDOfWzi0
iJW+4sKD4UhK0vs/3nwfOH3w09Zy4n2m71J81hJIhaig9NowTcCkkmB0zgTW8fPph/1LR+pJvXet
q0l68FOIZUyBjBxZPtf1yKWRUl5nSNgsWJEs7xBD9gJQkyqBKU3Z1WsRdjsIqOAIC0YqSBaJ4BUK
nV3ibc04jnvLiIi71hVoCJZakdyHiE31QFqbsCBmCG21xEWEnc7nukBQiblShrw9FOkAUbnUE+Pp
35oMswxH7UJrmRYxYlXKXSwX7MEZ4HSU5FdQbnu2ffPA65FUiPvpKvbi3U6OKXHo9Q0DDdXlE90Y
HNg3qv0tvq/A3b+zm32wTRwz/txfDypttRipcr/ES9Hgu4ueDkbRBKZSSjp03P+Skm9got4ib509
Z9edOMZXt6yD976Zpbk/cmCWLgMGgL/FBmTJBrwMrV80wSBa3uEp2zLAp15OKO9DaQaguhjZiHcp
XVvR+tlIib0I5+v23FWsMyWHvMJBDxeiywCd9OrQkpuo8Gq4O8YiMxrfOif2cRe157cArkP1nB8C
h1AeS0gumok9P6Ofp4X2V0TCg5Sx5TN9dqlxD8b4VxX40Z562KGEk0j83QkcEl2QnKkypl6ojVHd
Mdf7BpIXRl6nhACulCKGskfLhqP/AvnUeQZmAT9xLt47bp+nI4Lb6toYVijiEAUSOp7k+hE8rtgm
v/4waic2iyVfHrmyZKSf+/k1D4Ms92Cii/m98NFZD24MPP/8Y61m4ywPbMzoYvNeP6xtMlbZoRkw
msS1ynBHv188D1xJTGEL9tdDrks6RmHy6lxj3hNemceMngd/vWjm7whrQWFeh8p5xBwc+udzLagX
mMK/QQpkY3Ube32stDs1dNtd+I9yOE7nudw5oqaFQf0VQ/6epu2p90iGyyuz5zPUQcdzUCLLmm+A
ay9X5FpJyVYokIACwk9LWkIDZk20xFlCTD775qg1JuQVWAivvmPPxFQ5C0mvpoSzLmv5En5JUsSL
fRL+5y0qnv3mzX9sGkOFJ38ssJTdqRD4jAUIkYFojoBoU+rJyMFBmXhelqlcfBW91ujRxEMTxNsP
V87RuNcy72bmseKklP49RdW/MZ7lqoje0uY17z+s0WSaMELCNIvB24mcvk7cE8TnEPfVgsW8IWcE
rREqBsJ18p3WwAXuhg07FUps4r8+qE6cvmd1E1lgYlEKGAMGsime9/KulRWk1HIkurdqOgpi7k1R
zCGHqhd73V1kv2BRZ1hzq/NDLJFSaP1Qi/AjdVH9p7Hs33CBDAyqGLxphP+nafYIVPYfGC0/TtuB
Ij97MxGIr/DjRGnjLtLhTvnDaboRoAZWT9fSaNz3NwrTIw/2p0Bsfj14FsvJVWWD+5ENzTlypZdo
Fv+Yo7nnXPul23HnBDFhPkCgcARFNV2G15kDTCLBcF/9g/UZyAdN0jR/6JP5m8qNi7nBcX9UwgQF
bjifA0ky3lqyNcfmu0tKRv4plh58VpEimTVe6hG/ySDuVvMcWHN2Z48lG2tWe3V7E12qF3lcSCeX
kMcHoDX9XZkfwNanLGKXs0GOfra+1sFr3XprsBhjhJYut0mw3JYnmS6u1ohA0UpKzeG2fUeiXZgb
FAQYh5wbirzDz6GsYexNgslRRZJwP/ZU0TneCy0jwszFFlAPmXv/6ep5L9w0o8fIILhI9fN2z+ZY
8ES5ZyOCB/RY1GuJMPrUAokWYRkaBMF1VKagJx9QcT1OaHKW7uIZoaicg0ZmOxJfayt9/r3xLTWH
vSA2Gr/93ncMVc+F18PeMfzn0jXf6MONV6Ibeq/jGqnN5F1othUSpJkkTkH59mJEKNT6UvOvgam0
i+r6ZSAnneaLf4Y3GI6H/KVgY9KmrE4h0TzCv9Y6oquA2qjFHMao54wIH+1PoHJLEWmlUZbd3br4
rVHBhGeFtbjCLt0lCtTZ2xB3SzPmdlhwzwSJyzLTwUgWDbebEiR2++Per3sdHwlRtXzDrSRBd7rJ
1it6ggk59XiQ6fTpo4DjiYi4srhPKzxf42lZzy6jaFPkPw9gXpIFGIQYpDi7eIhVsGpaS4Y1bj7H
o1un6p8yMjbaW0du4O3JSnwHeM3Aa6olg3/MLGPj/CAYyjJVC5Bil+qPR5iVE9l36qIQibpdO58H
UP/4E/sGopXgqncN+3SOjeJbHbSwN2D3e1ax+XgPlM03P/VJ/GX3m9HfscQN8cJOnTxODfRJsfnB
8LYAFqtaZu3fUmuKPF0JOewEx6DTHz87kvlOhzQfukqzafZVy8ra03RpifhlEGhYgLiRdSddR8G8
Ux+55RQPe3KU8/oT35R8ub9FsGDqemO3Ohr52hO1LRQDL9E5rhtNraxUiyEojfz1ZCAcb5kigCu+
SubdbmHa7SHo0lB9VQRPurl+vwlE7Ns/cRK4TpSHAI43a16GeIhgx+8Zlu35icdhkM6QH4IKLdMn
TrFQVlxDS/4RTCbY71ooK35PIexZOYFy+KEp9ePDo5h2TqKPowFhA6SeZK7u5O1jMiidrkqzlCEB
/CXVOjUmE6Lur0XBSy04tJdlxS+QcpmWA0SssA1A9m8x62Ys4RN7hpwko2lDvLymAUvXzN+hJd0f
/IFOovxONf6TMvewsF/SPHRws5uuIVAeYSicXlL9BwL+VmbQYpfpgLb2lp4AlcRfbJH1aKKd2tf3
U81NXTnhpz3uDYWwdWWG4XrVGwNCcdsBVoG3er1sEtirQolFbltIPySXWzRZy1mGpq/mVxlit2Ei
cGZ9nV1L0WDI6lXK+X45DTqbpI3v91RDV3+cHNzYbdVOVUva8oWVAFrjkUYWta0PVrNIzVG6/1QB
xQPgKeA7vqRu296Esz1hfEQJu1XaGorrbfJV6SsNZZwF25Kvtex9V/kfj50/JR6Lf2ATjVaEjo1E
mfBrb6SFMPG3FGDfqdA1M8uEEqAw0Z7P6WZErEbuzyWIbBvKj4b7xF+/Egadopn57VnD+u6Fc3sk
1ttLC4I6WaZzvoacjWzm31A6POXMYzmuyXwlmQWD+7Izmc7ziI6thmTwZuruBIj3YntRwVxf8yHd
tPvbGXSEOods7Xx7i3cSuFB6OMGAO3h/bPqtdxYJDiFT5aomUp61ug5bY+7lVZFRvHcqXqqwHr21
XythPPtuljIcrYe2xvljoiRXZoTmBJtQNPFsrxvXDhUw7D3HR3e5FYbbzdh0m6qetHT+MUFRV+xA
LFx8tYw3zocNFvHqsjO/yUNFpCitGg/6DK42wbP4qRtiXPSq5aVEEUpZMGR+ENE1axBC9YA9GcdR
eiQ/J8ct4laPkDDdt1J6FgbWqK2a6XGipyiwqYCLTEkR95AlFl1r4w7NZ4BdKHiMgJBI1cD+cApK
6SHo1VCAlen6HsK3EXu+eFka5G5itO/4Z5n+nNCLWoI9m1zjtx96FL+iJzJl6BxjZL+8W3i5kM/1
2hBVIgP8opOwOuRn4JJ4ZmxnzMNHLFIwiQS7Mq/HajmZ+DZOxkkuR6K411/ddKR/QxcOGypitIvR
/z1tu0kKyLx+Fd2kK0yzIE7G7OL4TpDKJnrVzGx4VTPyguNQMljr9INjlpCdrCfp1cpcVSXUbXis
fbzn1rA+h1qCCw9r8ReqV1tR7B7a9qUIenRVKw9r41QPfEXopIwEUB5fMSeeSG8N4OKN8QTYYnix
2hFkIRoo9Le+Wn7Zxea0RQdR4UsY2VRTkIvPuu4tck6TmrXA4ccfq22D6KGxNZ7uM0GZJiquq9ik
TAM020Ya8iq8u434nWEPRuXRO7EGHkylXnQOP2MmCSZ6stEIh/XuRBhUGXWA0GcYCo7l4b6hHrY1
N8AzmGMWOVXMonIepzKQT0LxSzL7I6tmGpxV+xPzfqXbXlW4x7sksPJtfYTxM6EmYuVIeyJcsu46
gati0i1aA7QNOjImIzrpFrc+9rR9ZW0nuLOf0F+Wp4AFxJrZiivm51kNJX2gFB2qIQ/Xesb+nLOj
/YPInzyD8T2a7v1yNOl2s8tWnA5+O+eknzM4XFjm7T1CaFN5ajqfkFRlOsN1XsQ5RFkgYfUZM3Pq
FEBZ5st88gfgXjZ3A82kKtXveUbDgBd3Q+fdsczBLRCs4qZ1a8i9lAN4T5+vVoPZGdzEWm9wVo13
IEMjBTzveaK+rgRXdjqUXppNah3HWLR4FCYFutPumTrpdz1T9xeum+S70n04b6gRRyUxriP/lVqO
ULWG8bWGSKK08yGIQgd4BMunDmkR9R0tAws4mtqDS2IlJ1jiiHxt51m0vHEutgyCT9YhhUWkcBNU
PDlmuWl0jEL9D5XdD4vRF/VYnjBM+gWMgsDp3YUM15CxucV1Wn4rKhv0W2DYDhM9o0k8hymQ2E6d
C1JEybvpn76sTqsjHL8WtH6GhjIho+xalXR+gaZDEYGbWTzJCdaty/LMXaQUK7GW1R+5UJmD2UXB
jrjpC76051yQTrER//upXhfI8tV3aJuGilI1VkBSXGpjszWtyA+OHbf/EEAV9qNfmeeaeedS8tcB
XlzobBKuh0o9bmuNRZwguxs56hyB4xAGjCHrnStxfTuHjLoQYY6Y6E6mdNvEayxQJVNJjy4Yj/rY
hio+cc/b4+GdcCnMuiU+Ikq23ia5ZD5L8JS2vosz+NBe5JoTURC08exZMi2T77wH2Csfl3DJ7ajB
NnYgIz3mEaXhy/oWUEnHC2hDHvJVW9q+8+ibzBeoJ5zh822HT0s+lNIiI60txGEQ/F8vrETymHvW
MNKFBogWTAO8kpt8c3KAWslisphw9UGajIdU9PjyDM9KLmATwwWM4uBZhyOmvGb4GfPe8mdGqQfu
Vvx/0VP6ioMf5+Jb2Eg1BclPzc8TV52WIne3qeAspcSA/o+tL0+K8/DA9/ObajZXH5kv/4wO1iC6
Ce+5lAPhFoKZ5M7AGt7JbVrqegFknQDW5Y53sy45JjKxmwZiWDXALWApY7wgItuLefVvBySzil3V
jFrg9d92HpRyaRZF8N/enEhAaMle4Q+20tn9Luc5XAy8ouxgQz54kxDhA1nbpfn673t9+OfGs19d
817g/MfpcM58nT9/EQJh0W1RilSOL62MIYuw83ebrOCU/XUf2SUA8/wa0PHcnz8SQ0Yj52Q1dH8I
r5jsKZASyGK+GdWdtzkWUAH9w+6O43j7qVs45S0qyQpYlGTxDf8Vj/hWR5crobFM8oNLic66rpF5
fltihHvghSA5USyt7AouS78peSFKUTbji0E13qQh+I0C3Wimiw/1rMVyexW/E5PyOWxGC1AIV9Ss
WIEspqrXWyBeQrwefu3aVV82bcc/LOoEGHKeO52XF0e4gLdDvPKKEwB8muEnRQ9TBtNWidQqtzeo
zEFc99kLMBWWJ2oZnoJoVxPtVa22fG8vyvk6DuFmV38bY/tuf7ZoORV8JXoqgaPVKGIFaZ+RqEdf
ocZcFto73RIZlOMKsCnz9P2beo046lMDFiYvjoAVsCakAIDg4WAYzsmtnwMnLihVMrlBR+OSDWqZ
QtJPxkkuX7wJ7kYs+hv13W3Ri9EB/OrRp3GAnNPGP+vMQKDQEiJ4vghsJGhI4+vcWGFzgDuy5zcW
lyJTEDnj6+RTf0T0tlFvSWkPRcuRc9L5AFZLrL/t6NG0sIolv3hv3GZ01PBtuSGPyqxcBrKBsSXL
IgCOm0uxyifDrjXEiV2pBPsR6vfvZKHfaD+4MmjU5VEvy6iT3K0TeszIL2tp3SeN7iTdRWK4hl6H
mQZj05bjxdv3UNgNz3h/aMW2UNHCEtSJ4uoUGJcyg6YSY5EIktQh4jtfQYLVOnwGKzOtZVRJFoGH
2/+1PGn4IDn19gQgJXxAff7LgtxsHwyo4gIIf3366jlLTZ8IddNqhWlprxyogjojHKmNAicgjyA6
O6d1LnCx3/Q1K6TFzB4BWYfQwKiUkWOIZrzFLQ83XyMwXAH+yq6oLbx4+ajZIV6o/6ORhiwYBGAA
CW9rWh6pmsdzUBmgXXRUNeCnoj51IrFTNIvWIE6+LIQOiBt2BldDm+wGsQbyUqWg4hkdqxUHiFOI
1OGFZf6lAO6Urj6rnOCIE9oLQIGrs0GEuLCs2G/Ly/UUa4AZv8S7FNyML6zQclCNbphz3YS9UYTq
om6REdJr93tSu3GYWIzJZ6fT9/WRkki7lPDh1NA4rlaKntpQ/yXPHT12b2kSVYR5m298yYGoL6uN
dEpLaP7DfuaR+fvzJ5S808kbUmQhB31IzRUr49bl+uZdV2c5KEoAVPiCRl1l3R2Kwiw4RcCotuj/
KxRmE5afUCzaejSb2Z6OHtuNwuHKp3JWhijyFFSQGHMTcJ+eqyTtIAgOKfe2ZJkKI0dzHQ83k9yL
MiiIGgjp4tvxQluiDEdBIIgTJ/78wVG28xKrufvvv7egBHC4AVowjU3e7O3JDTseW5mg1o6HRmau
Bvq1ClXYkCd85zBWO6lDiVriUgdJw7twpEN77/10ozf97BRKZGKQ3MvmdBV1QHLcirtHvuTI8DcD
HAly18KVjy4l9GibLQiMHNJcrHzwbe0SSlfQ9Y9302XJ6hzqyR2lN0LGkwn/7SVvpsZSNpM+w67R
2iFvmVHMQ7MmTyNBdZriPcN6alw6wUaRzUe6RuCfFnUaM6T0Z7LqFgGITGrnnk0hGYGwq8TGKAkr
BeLH2+HJSLowyYNSRqcrClAxcnqSRGU63AnvSj1NMi2eFXN4Wfysd2+QS2O/JGCkrZshh7XvIIQn
3JaVmTjDWbpRFF1Dabl4wT25mLTOT4fq06H66XJnOIqYgZYczO+az63wsB65XetOqv4/z/WjNkOj
5wzwTkxK0r7+0A/qcOHtrnOrxfrHg/UjgFc+dANJuYG1NQwy5BFrhxwkWVf8nXrmg5OES3Ipo8f6
WTsKZws9ki3KNkg0fS8fm6XUVBGodicxiofi+N5yq2YQBCWcI5BAnD2AlfSlGMUDHzsJVeew+vXM
/8jsdnpUkO77onRz4dIdRitJLkYnIYfs+mZxVicHGBqFPWOeyWVPbgsppdtmI/jz0G22OeiRYf9y
1vfHNWhYdLZ8xbzZrHmU9f08hYCRsQNgSrugNdrp5cUF7jhEZBR/yTT475iS5uNWUshbHX4ib+Fp
gafX3Ip3hPFTVJht2ajh3+fLoFuIlioxO2fXiG/wfGSfBKypUoTaYYTBUlROqgOrSzV28sk6Lw/L
KOo2kxDMPATzRsgkKfj1H/Tp2MDzgVswWR1oqP3SJfJNL2eAjJeZ7q5HtB2xuRP+GZoal8n/aeBW
VNE5ApomLvxntXwW76EtlqsuXJe+CzxjqMUXpdJBY6Bdlrgvsksmkq/XVWcTAP7omTMcekhT8ult
/re9PaAYJnttOs44lQXuoM39pechXryv00HTq3JPiFKqnfhc+pxQ6vwdpwEbN6GHLGaWGyGIHZpb
pc6/jTU73O49Xme6dF8W4TCcK3ixkZdIIVsqb/ntQ8+wPztXK7DbKzcM76++gWzv3gqYXTgFdFv+
I/vhO4O1Gp14RRXtG85zpxpFJs6iWjuQiaM0Ce0RJKotDNwYOPOuSwoIolK19boDTA4ZUAEru3SV
h8avlx9671wpQtngLUHCR57fwSLOxpz9zESgUf54ZZHjW6zEVrzhTqe1kmsBqYGBEeW164y5T11Q
gxzqjApUoShW4R9D0LIao9ozW+3/fDK417bbcP47Tmj+Invfrf1c+tIKE10lJ9m81dyw5h0l0pOE
20D586tGLCZeJaJ8J9pyI+034ecZ6CI0vk43uQ8GR+jC/BxCVd6Wdq0w/OUkMv32REYiLzGxe9D3
k/WUYbKZY9isZ5Afbf3ArxwHvwxLjDyceF+ZCZRaCrd7uqNqzgTUrsZMOPANh98LJ8pjOFUkW9Xa
pWH9QXgNaoYUDHv7QX52l+uTQSuotyZ41vIHO38dD1+l5gMV+MYYLpUwn2FDHNgXbvtLHsF6GkfM
BVKCite/TNc3V6mIIFVOiJLynFHFUVWZeDzQyqtxDOI0wVW7uCPZNr3rZmKq9lDA6LBEydTvsxZa
UGUNUP4N37H7ASCWNouFPk27gjY1GPsCDvI/PsDVoTHhqAQxWAr9FhV1y08a9wNMhgr4j9rGSS7/
aal+3SRHnyoyHJ6KtyQ+/2Fa5n15FBGFAtDkH4mDW8Ie8nlEQPMKhoNTfT4yngxZeMrqxb0V5r0p
WRuhTDC7ZekayM6Sx4VT3ik8QkL/xKSHUYVELscwdPcCGMjPHvHDUV0IRgcKGChJPxGAN2NxAIJy
6BQY0Stn+446DyEyae7cewTSDHIPPoAy2VvZLWL8IXDvayRuspePSP8+SxOu02y7f2BG6Ep98jfe
lZrdXGPAMGUXU0ZpJoinTCB/f/8iy0zx3gEo6AW5FtF5MgdHeRLZGzXxcO7XZyqPFAKKK1iuMZ8D
ROKRoBzLEMPX3LBxf1fWk+LbUz0/i0xPCUJSBQsZy5h/hhUcN2uSMvhVe5yjtDQWrsH9Au5/yPVU
yMPuOCoIe7cXfFVtxN/GxRzjFdaIwH79+AggAQ/Q9l4NWQCkjQUcGtSwVNO921lG9yLzXGTzlG2A
tdQghfqWTaYz73QkQegHuF7ZvqZSGYYob975lIS7oFc6x0noVzKJmgSUQLNR4dfREST6Dv437H16
rhfQGNqoji8KRcB68PL2tTlGlUGKQJCu4XfYxjZfF62o+8eChhQmMAMNytQ+1s1tfYB/6RzJvqNk
NZTxa0sX5q7B6EO+ALCob4KHNYRJhEqzknfLiyMtucjgZYxgXoMEtRrokTcEe5k+HZleQwU8pQNK
z8y9co3ex5C2W4wkijiEnHnfghLSKt7e1PPu2HoTZAzMgLk5vvE0b5NM9qom519wjBJwzpdKN0AA
VhNzU+uzMSKNKqkMaj5rGLiAKpnNl6boAe4N3oYI6GE8f9EGijRmj8kIPTjgmIsgzPpDVluX8GQn
pU8ZzngJ2pQ5sbMv1l8lSSqO0SnKu+hWMr9klhmWbvVgIQc1b+s4uzsNcdDq1L6Uwu/6anX/X1z/
pFtNu9p/NLCW26uid90yHILYTw5a7Jfzq1dOoWXFRmtKurZEOlknpyyAUN8UVJ0VFZN7Mhs4yayU
jcVM6cIFeskBdGLCrBGUgUrGlVOOQzvNaNj0mN40Z/pdYUu6FjSFd/2gEf8uq2YqzElR0DmolMMt
jDy8hYxl9bD7Fg33bZYjukV4EirbDXLnGNFeOTVUwxXudb9tOEGeB2HfIinKSeOjLdW64hnz0ric
czsSikHWaxD9kEh/w5oBceomk7q/14nV/PmJNk/hL2nILzTqzlSAkCaLO29M3Hds1EharLOv2pFm
MyvQXvOL6ebbKBTyeS4asz+lJnj4PJIN7s+7n5KdHUslhwm35gZQlKjPOF4jfPjxSYbefcwTFqFN
wbq8d+kXqomnFZuYp6rYlV4g8VK63RR00iJyr2mB+A3zNFmB15RLnUeSZVTp/hkekx/jg2Wk44HB
e3AVclFwRkTD90jIW6aiUm/IO4HBSzLJwciJK9+zOUgrioKRrVDvzoJfwBkTH/LJUbCfOSVQQlDG
Yx8qMsOmCFOVomIOJatbkHosNOGaGPIUToIJfb49RH2RH9vHEQJ18f/JBy1HlIpU7zOEY7HEXbrH
6pQAAxkQtGrCJB048digSIVQ8/GO00WHbesvq/62dObc5s/mX0lPZ16s3FyFF/GCvCEZYuvGZVsl
UoljZYIf3ZDJMjgwvlZv+8carUyOw2Bibz21fV8QGtiox4AnV+4LwO2ek53kyFUo02hLI+ZSjLJo
/JtuSXlFYUGgGpZpI6fF+QCs847G1LrDGQ5kLryMQiCWIQRvJzGtPr2Vrkctp21axcwl9TXfUapP
qKG3/kpNkaD3pXQ2eHViS4gjic05Uo+FvOfV6R3QegPGFKFF/0enimTu0NCDvjjIXNijClNhBncV
rLLOf9HpeIE/HP0PkrFiqPXIpy2GaluXk5yZEtYNcDOWtD1PIqVXT8vO21sHP0TllDjb4cPWCSeO
+uACJUjqoFHzQyAT3iAHEsauavOXyacsA05+e1qX39x8HkvYKGTKjtLSBIaQlFF1+pqMK1Rc56Ay
0dHqjFMDgbkQlIrH5g5zti9KwE36yk8+cFhNfu/NeU9eCC6TUbZpn4iczam3mgxfcjPucr+6m6be
2g20TIr2ExN+0MunAKYhjeAW2+fTcNbSYa24WzrlW5ua9qWFCTSTFVq523+XMwTNwc6OfDIQ8aXj
caCpSheZzoFhdTVeGpIC7vqUuHqUz51nUbWrBkIwG32RKAsxeo7icWmoHjbz5hhf2dnRVnIjd3YW
5iS3nj4J1RUoQk7ZiPy0T52nF1r+vfobosyazmXybo9Lgk2lIsHAY4RRnYT3XJlVQAsbR9/4CaLF
r9cOizL9xxQv/Qnt6dMFwUmjbNmoLkZKImg3UNtJ1H4RvrMbCkeAjUPB1WZKFhv2CSzSae1ttwPP
GD5SUwGoqArVHSsuQc1dO44btGP4esty4Kloa0CJY8WfJrTeEFb+l+M2Dk6JCfHvA2hG+3UQAelx
weQAvQ12R20uB3vIoZMwbRIO+h4+35WR47/NVST9UTBzIyZlSe4usxXkG0jZlgzR6tHWn2c2pLVD
5/t17Tb6TwWgTPfX0XWPNo+4NLYwwywQV0piFLo0I/0n449bBNxYHwRTI/mbXntIxT+gTJAjwO79
ogRjOu0hpA0BugeI9fVp8ddSOezLL4xDF0PcXyi+Hp+PeJCpSQYJyqIMsp9/S50SmxxVa3ytAxMQ
ghDpx3h9kOWmce8AYPi1Dp6dF1dbhGWXbrzzCYCGQnLVhqt+WcuOzWzI/LdXNaJedufU0YFT2tAO
NgVKqcnWfaLlzQg+GwIvWSe7G3Il7LTcFIj2usbup6MySLSTMWYAryfwwXvjRQMUi4B+YEL6I4Ra
LREAmB7Hk26buAJHjJ5m7KeCi6NeRruBV6Cv3xttCuFklqrFOvIzU5vVrHgkdwy+eXKt0zaDpIir
vfjsviyHDPDSp+pDv6h0alL3knYo/IHFmSM/jieJTD2EPSEDKY3xMvqrIYSg7frqHemOp2dEthTS
JD8/TMPJelwAbxCfHcQ4OJHHfNhvSPgdHRTP/f1vfvpGEQ0nNSvgNPYuSiZs+0IgfV6pD7No2kWZ
RWsm63GdXaVItDqcjq/4rwss557bYVjTZaNG6jiOrLD25aHEWKKJ5sdsqNwfthvZkSBefExJ/ACQ
soHK+CGQ2iTzq4KopAxHPowd53AP1eEm7bPEKVCtaAszSSVFbar6SCsQmpbM7YqAoomgFaCc63gd
LcViB7ksRqfuf5uUWw1Xx7n516jBRgU5f9c7svW7QKIrooNslks6SbzDQGvfFD1q7sDGJmej6Rjq
+qRLuuypg/qWm1Hog0gLC3++tE2NCMedYMa17sF0jAWoDBUtHKkHteA5aEFSlaKzOGssjPclkh8h
jawdCTaQ2T4k5yNvdlSXh0usyWtXbcvC56Ux21LboC8sWgXdukd6RWni26wP+sEUhs0YfN3bUqwj
l8wKNSekKiE1N7gfAJ6lnbs4pgB6vF6a0xwDWsNLQDMCerhnRrhGh6yVv0OYJbehkwMdSjsOVr3O
LMi+1AaftoUSREKYRIC04UCq9o7CP53Ty4l3Xp4ijT9mx7jEJaJnu+14UWVWrQ08T0ughLHpDRF1
1VfhGA9uH+n1rVvmRA7097LAYkemM1GGeXlpx4DKreqE2WNGpSZ/X2BHuY1mldpk2AfbfliTWkHV
G6OCiCRnBA0gjF+yPVXjvGvUleO6quPFWPk+3HuafLva7nudnFJARM1X0c5x6bOe6mCog0E4iubg
JeOU+5h38qGEjuyay1lIBTkT6hR1EVn0ImXT45DVAnknmTOAUL72pCYfS2KSGNnSo3Z3AOxfYaTP
7+1V60BJ2Yd18N/FwVDrtiUgw+Ujv1wNosUx39h77fHNHdU+n9MFK7m31WyBDQ3vJmwjalCZTKzb
wRHcNb1QZvVRZLn7trQeznLer6WFi+zGtLg1OOG2MDnqrco1+6u5cjwJdsfXBVUSekt0mSF4h+oH
L3YQY37tNeL6lipDODbHoeIehqfiGSsrxqhxQgSGDcLEBSt4nIZbetzkP37FRZLYMcCEBPDQQsmo
VtiuRqhUNd6xvQ04FUiYX/BntL/ypiYOnPEKwzJvr8NScPqCKcJK5fXGfP1IYyNrWtz43Ep6IT8k
lYyVRnzO0i/GIApt4m1UWnin/7XFvRyVpAKGITtcpMnETdCke3TfJxnDDXp5cmjxVhxqp6S4CqZt
O+MSe3LDzxmtbjQ3xTQKxUfRzqu/QGFeLc5GuBu2f8O4G0uOJdiqHNibv1aeT5Bzj9F3wSRtb+r2
S6UsO2lfewtNPqrnPSNGYq/v/aqLWmkKzeWX+zPpFbOY7l+RhdNaWPzDzTmwXlaeNvhbSJsA8HkX
HWJeRtuyYXIoFHRnNOh0vzqv1l4lMnDQNChzI5Q2JrpuKbRHB4vwmDU6YqEu1Ox1oDfIashL3rZO
SEIVtVP2pQpqBmVxQVKiSemt66xMSjXLYJ1FF18eweRwYvcT8t3s5y5WYzWWgPVo5PGRVvDIhFww
80gsuJ6HHiM6sWBZ3lz+LvigrrupuQiVgFbgKE937JPEm6wmR+GhB0/Wk8N7VZEaTsdLLJ9TJcXH
4W+tynu7likSy0mav/4+7WrTKAlXxt9PMIcE4eUASLFug5Vz+JEE6fsNo3d5Z8RS7NCCNP+QKau9
FSuQRI8geVtF78aQ72ETGWPKPHG6EBIM4hVClpC1A+ig9LdlAVarPnr1N64vwAILJqOo8xsHRc61
pwe4wKMMdREweKrJ/oeAoM2ir4Ned3LaQRhwQrtNYgqggKIpHKqtwruseqEvBWJmSSfGMw0H7LdO
BeEcbm/Eql+pxyioOOMUnUc0txzMu2I2INYVAHbrxivObPZM1zCM6r9bHvgozEZsNzN3OQRQqZdE
9ANx8tNZfu8gzjq/fxq85wgumT0YF5uCdhDq6BXsRXdW7AoDVG9x/XvC65DR9knSP0ZJQ0ClLfDt
SIb7+PdmugcTgeo0TjysTKyP/tu1JwybkbLotKXyL84n5UDxY0RBoJ+MhDv117e4AbXhyTthoAiX
1JZfVtTrWbnA5oovrKBEYyp2/YNBF/2bATiRGYU4z3kBOKBRGWqFpEgiP5Pmuv4k35xlAZxef+hN
0H/c4Gw6sOjEVqc35r3GuRTm+dUZEFSDhb2Wgfz8s07J9rSyUa0tttH0Xm04HDAJhRJ2hlfvPBHM
9de8UxD1mJrWaoL/awIqRWi/wSbWNKz6EdEQUn+zu9MEwzjFBGteGJpWqy1hsO8YCd32c9RiOryE
fd3UX1NipsycqPtu1X15Nn398YS/pi2TmEkwCBFxRQxrCfL6CH70xJf37pSS3f/26J/7DKKjO66h
GFgd0LB3SczQgRoZc3sSm31kbmD0cpAoWoTCVueMxddUCLOhCNaYyN6xZjIApzXCKITXkCjDeWsi
xRyuS6GQNwFmfUrQ5J3mGFMswDCDh/ngJUF6vWlDD+bOoz85AjYGPmvb+axzz6MPADyug95OS3Cu
ldJ4Ln/DDosbEM6x1G7DdmLZqZpVXXpHsVSsqlelU4siOQ8zXpeSpnFbKftsWDPLpunddUPkPymd
3DxcSZ6F528yV/ye8hqCDnr3RlKDldFSGNxmh8LsX9yzYMG+ru/a0zFaFa+pJmxBb4JacLJ4aFNF
eqtxoQk3XkJ4utI6Y7a+/sHTnxscmcty9ETfE/zkSckDKuPdeJzk9BlOhzObXyuEK5DFgNTN/gSl
DKW5HHwmnq+5sRQhwXgNc5RtUTMgr3eyx+qrtyT1hbeyZN6lgENXkTwoGXQXiRhD73zNbRDZ38Cg
ORVu3TV3bDqViaionuBGTx1typrpnS1C0Yw6CQ9wYFt382HuiOjz7uZtGeQziVPpkcpTVLDREi6K
jqy1bKfRp1CWuDIJfKIGX3Kv4eLGEyd00WDBSSM9c9hm6EHW4mC6/SCB56p+AJ8r2TZsIxfEjEqb
IlnutNDAkLPnAQKRGqs4WRnDt0yXcd/JpPqi5stWyFa0P6wjLFRwv3wUgoFYTO281VYNfDMlKJIT
JaFjlsxkQHP/sKrTuW1pY2dVQdjQxyK2F/IAT3vfDLs3/sbKi9kdR7Gpx3gbpi8KAi3fQ6nMkcxO
+h09VutUpkGJdlVzjbbEcfiIn3I0UMFKHTV1azUJ//w380aOVDaXRnPx624RFKOCHSAKFL3Kp+Gp
pz/9ckBYVPXHbvOy9BvYz44pkF3O/d7oaCfGwrT28vg3JTfcuz1W8G5fAulMwNvsZV9cJJ4qWdL0
3e/SC3w/Awo5ytAfYTJoOPtbHK4x3F3Pfb5XJz1T4DjsHMy3WYU+RD1XhRnP/rVZZ8GFdLzXlfqX
fimWbWPve/VOMHsvyr5ApNEoOQJgWbwdPGuENwctO/tbIxly8fu4xfzEV7S9kxTINsWhLKcJNcXr
KE3PFAaZci/pdZ/Kp8QP0o3ZEU5LELHQkMdah+BWziFYKOCjvK1ePDs0wY2ygB55j8+Jcg104JOL
D28Ya1KC6G+Ys66WKuYVFvdImwHSxwAwxAbN1D6cbQjnnYyyOD4EXiJA9AQhfaS5g6S3Ljr8hDc5
VeP+UemqLk/dNFxCYgFtPZ5Ytvo9QCGGM8RXyRA2pSRaYalYSklUbZenZkmNOD88xAgHAof/cM2a
exk0NL7k9aPLbKXHgTXtodJ9QUY0OLbLRTJSG+3R1XwROgg2Eq3WsaVOUVJ0Zx4sIaZPS4Kylp8B
+IPImSANRvtzTHxBKCKthep2895xXC6CyUM93xlwog9QNIr3C5wSjyb2NOH7eNHs5W71m7lm/ulH
Yzg7rZxoUSOe+LPAMDZNRrbuL4FNKi8C2go3MNNktBHWWsWzvfiIpLNmu+Faj4RkKiOtdNCgnjSt
RHr4QMiZ4xgXh6DPWUbxmIw4akyOwv7TTmMHE4WGv37klJBMl0I2s+cup3RaUWiJ7ivQepPGmYw3
ALD/RLCmOfem+VBUgMRay1FUBscxnIW9VdoBOHQRegiWkqket/nMWMIO9JIr1YUNdmc+WdYaC/ut
k+C1ptjxvpLJ9PLDZ5PM/O/eBlSrzj+5sbAHm1Yc1GGEnaL4I/zu9gsi7Q9/ZxJRKpSbvlDONqXQ
zbWdstH6eSLpboDHAKgvK3JxdrGJkebEvimE9Q4UPPIZrhg2YHNoTgN19+Z9nqTholfYDxqKULR/
Y1LWW10IJLlFv5t1Pw1eFWeLpMtzKdR1yM9hV6+sW/2GIKL8e5YRjXKBZzZDKhT9PUhbZWGApHoM
qA4grOWSzt1gepPuEh2s6oonhWzHdpsxtcfM97fVfOldSR/RuZOK+1NxsjOR7EVOFoXJbgMYw2dK
72kW5jQsjsarNL0l87bUhCppagBxt1RxLu8HjBNBfMT/w2LJiZQnK5USc6mo+X/HIEALaylmzJvD
5RLaiiLKbZNGtTWwBJ0qMeopwxKknrSbz5gKCnELJKpSulO2EDmNYHYbRJV4Opr0sSQPh0CijPeD
tjVtiRHlRkUHCm+v//LGPPphBSY/9nmCp8oupK0jkAVdfJkH2Va54Ivyiui9yS37Mn1INZPJ6q2n
N33mFHOwLVndMWi4u0ThBrw6yIKaauyk7igu2RclOrB6w+n7HRtkBgMv94mwJBDDk8h5wrzwjCM7
h7f9usa0ZMJGShCntXhDhoZhGKp7Luk1xis18+vuHqN/4Frv3TEt41WO7VX7UFStKUV+gDS5U+7B
CUDG4i71BHbj/T1LnDdImfHxPkig/f+W+jdiI7dawDmKjUQ70pTgfMNcYzP4Sd6dyZCyDhwwbXE5
Nf4H0baAH7YsLxOca99ArcMnUitaX+DlDBCaT94Yhpm5ps5Id2BTPGu/kWG1Ik/dL/JZDCpAclkT
MUh/8aFvs9jwunlt3ZEVzjnXqlUyy3VAoquwJEpNCQb6zrSPhkuXUfNTDLurztrLamBbwibzLA/G
/kpVoZgGLaZKtxpzXhZ67oseE5LFdFD/6ZDSJLubkcohCojaMx6Kx93mAslEEuF+egzNow1tNXVS
O3bXAbXXrq5gRA1fZ13FjF3VDvQUE+/p6NCBmWCKpHL9B+W5XLlJKvLRiKqJyW42pNujREDaxsYV
NL+xrmdy4UuZ+rf7eK69Mh88yp22qTf+1NFMIboG7nC9dWsMd+QUX6GWOLrHaA0pxWEUUaG+0Pg8
CfoeRe4Y64+v7ha2zxsBFdBN4TaDvl7EqU4C7VItdX9FWeux2xxj9BpSmuiKy2OuK3Ay155bTW4V
ysdQvwQTJdfho0gCmER+hE9FDdjp/ce9kLASvCIY9xpjiUkgXDiOGVavA/qc+2GkvEUvB7g3JN5M
jrn6jEaJzCBRqXC+fADQpTNj/pu772605+8FeF809jFBHdOe0tjrTLHvD/Pd3WjCxb0y7rIhIbST
lqA0tRuCWcNuCulpUsb8UDcgXlcNU8lWGYUZkHm+hrI/mfJ3G/KVz62VSrNY5NNqp9m1GFiDtv9T
Po9T9Qd32SiCr6SGnNGdb6snfUfqo45+pLK8oWYysmu4Cqnjc31PdLJEDRU2lYJo1ODGJlNiiE6T
q96JoXQwCtXK8RQ3KRI+quJRetLIEaRQ4OtPW4jhFfLTwcQEsNiD8j/GFswAnTVZjU1VK6Aw97xk
D08mr5ia1bolBK0YE6HWBckyMbtiN9faVKYHB2uEmo7LND59/oj5Ind0y3mhVP3mdYJebElrtrfp
dkhSNwy5HEtrVuP8F7613Zmp5tWXykkxiloVKidOHSgW000dYa8ACkSs1gaTOb9oDdv01UGaloqn
9a21T3sEXhL+ukcaoyR7OXjp8zDywuOTVJKRF/EJsT83IGwULZ3u7RXypP4VQPDjndg74xqNqsMa
b3R9bR4d8J68mWWBahwfT8P7OsErWr6JluTeY/Nqe/SVGtHgskmLpMDRUDRuhSbRXNlIiocdNp9Q
iU0dzxMsGyUBkM0Q34YXgJG0ADOJvxW5iuuYEG7Chpq1vbBsMrUM9AfViVGfpWiDsJ7PRZnoVy0e
k2UGukXd6Yx36DpceBG8TVtvdk94nNwN5DeDzAq4IM9JoD1GVWRBNCWhmqbwBIniKdutEhsPg/jT
rXKhbeGtxr2pvrpaevKNz4Oggg3ggeN5Dl2K95M5B6DZHHwPPKi0fnQHmVJOj7P2zVbOUVQ91Xad
lqt7/sULUyEi+rzYMnjtt9tAaK94sxn0oYYiyvqpj2aiNUJUa5euc2a+/BVLCO1mRhvB/xxpe+nI
M42/ZbhUWvZkO+/54B25hih1Han+qedAIE0bPaHF6uxondzvBfvT7YnNucCiD07CxFFCyF5LAJuG
9RV0KPADJ4XKNHSaArdoZv4GccBBrTAgKWamsesRTE+L3eYTbd7OWtHiOqrwLoPjbummv9fiI/M0
412N1aDcNwWiXkEsoUkiST6RfvsZdWKwFh1LhtNJy9pKxJvT9BXzPzU9xF2mkaAMTrvckNyVtmAt
ThgMGcAOPBe7RCQdwJ4wF/UCrr/RJVGVU3JcWpK8T29Db4v5f3QeQLYcqytmuVeXKVJA2ElVL6qV
J5gC0ElLLQgk34dHyDl11cCQByFXqvrdJOYnDhyJ7deXup4NUFMFWWOVjksFmvJDABu4MFcMCYH9
NEvKVT8/PD5jSMh/gLSLc38shpYtpjLxpf5f80bjzTR2pjYEpcqv9BdkKwDpss+b46nnGWVsj3n7
ZLKs/JM+MddOTFkK1MPJqJotsDMmYg++ALKMAklmujyNnMGgxa02Rtb5C/3Njz2C1zxM2kXz3jnK
djmqzBhj8/WfJVHfnC1KJLo1runMi0VJveT8jb7vdHchYlP5N5yZrslcnjBPDGTMK8HXaVRDNJ7B
OSOeNMskjImZxZLDtj3GSa2AwWc7i1uAHxJlHLWGl1OvCoxVMnW2vfxO/cTBgNE/NaBWzZL/CfAR
2NCP1GJir20u0DkXxyQjjxGzgtv5qDHwJKfihBCqNe4LxYUwvF1rq4f8IWxGf2SjARPVh5KKL5Ws
A+tX3TaB3/65c8OYj/2mD1/WGOzdTGuFaOHzsJlN4RneQDs/VUGG689B0mO59nLgZw4MUg5F2coQ
5QjkxbkYOSZ2UC+qG5RB1YLE3HEmxLaJgSComRoopo2JLwPp9liW+vQV3VPmP4xSSFmM5BuOEVwd
8JQuJ05Cc0OK2N6D7nqkOkOseeWChw9BGVzEfDB53NbaK7s7QzP+6IV6GTrIpWpM7BexTGaf8SqZ
5eu91KfC2LCJznqw1m0b5Pt7LOWHiTPSYsTlWQibZ4uiID3X5ji6js2IxzFoF35JsdWx1eUo9WkJ
d4sGcxLQH0tIuiIpR0Mk0sosPouwc69IAfiWdZBXfwl2HaiCr9ZMjS3i3owIOIsJDtnb3Dex7u2G
McROomMSi7t6zX2G5LS5hnLrpK4k4Ym3GhqRXy65QzSJU1pW0dBiWUua1SPRWER0FzF+gQ8oxbGp
GY0Ahg5eRlkbUQU5uCJWL0m3dt8AFnwkdkU8Igm2IqpxfG7ZitHySrtootaMBfs4KHTJxwG+Ns3a
9reS8xFNlW2CmyhUrYl1QPXgsLm92amJp34dg7Z3XDuJL267YvS3pbA4vDfey/77nDY7BsL4mflM
z8Rwa6E4D8RGvgoMeo2MavEuwI7l1tD29pAEsVqYKAIWW8+GxwSj1AupSQFp1iD4P0vxooiqicIv
j966voM7njdYkRMCuZzlg9MSLbZYEs8TOz37yU8zSbjSXIPflcv/aF0ewVAHQNA7wYEx1P4r+sa2
BZ1aW40NsXkC3ZPtTge1O26UeoC/pEYcrqFjylI0LyuHeoJOLM30P/FV3vUa8+6bGhAermsRZXiS
f2W5M/Fi+3mu2EDttF9RuPM3NQ+jGFG9WSnzIzODo8mpSYPIq0zQk4rFfCQ9CMpNVoqQQVAgNKnA
UtsdXJtCiHpBiUgsN6PpwnuEJdRqmr2oQ9l0attmJel/ucgz6MoNJA+Nhj2YxBoCRU0tF9u/Kun7
L4dp/JDCbF6wT3qD+Pbz9hYqCO3T6bcuE9dknBrTTDynfLG3P+HmLyBUF/FA4KVN9+1IKo3ZOAH2
qmxo8hRgS35tlbiPFsP2A1v/PpTa/6HAHbuwEiuWWjy1Gu5V9/zVkjaq4wi6ZmTNNrj+Gr5iPdNH
YexPz2HNYWiHivz9HIbZUzqjk0sqipVQ0l9WJa8tEDg18tsdi4svASQcX97IDg4d6Vtil+mUnpei
3jX2klPxKhGXIbdEvFCUaFTTer+2zpklvgGBIg/rJUHWVtZUvlaASeqVDR0pACEroyKsNIcc1sX0
9VIkXdcCIjTpQmmbfuKqSMdWPdKhEZKtvImn7l3h9o847sgvAvAslg4qe7SfyArsTKZTIhA+qeUl
Mxga24R572uIA9HrXwIkSn4R1C3/cDhTckxFFO82vkNVvc/TZo894ir8GGg11nN07LduHxM/zvIe
bZjBGKfdJy90H8xHJKsUBfPgO+tYXzBmjU9RBFs0QlezwtPJFabaP/OAyfLEELEBUO5s+QpS9uMC
cEmvKp8HhzHiv3uwKcudFoPNhVD7V3OTGiygwDDFxUqNWC2+jsnB91myCLTSqizHTgRzxsWJ36EM
mCRDiCaEFTjuAXgOm0JAFdsWxS7LvV8ROKBEDafWXh4zatza5Ha97iI9VTYvK5r1LnQEe36fBGOJ
hVI7pJ9BmddO/a2aCM+sU88vens8qqmitDedObDdw7udUU1Q/beEoKeVfnyl5PaBbmQFCqDabfT6
c9TSDiY40pWmq4LXTDLDl7nt863RoJ70X8UCrmM2cSne3nr1lvAFudL/x5T2vBKnO+pD1/fU8tsO
Iq76jnqR64kcIRbmML4t7RV2aMRdwz451HK6yzUvkGn5tvuOnx9MDzCR1G51Qp5SsA+yJ+8/U6U8
3eX+1+Qp0sGOgzU0xfOC8POXdYZpT5gr2+XQtz4fgatbka7S8XYyoBZCrnbmooLBm5EsotyITIKz
Pw+qrbabqmQl1XEXvS0164fP2NL7F+1U+c/6sMZvh6TS+5c2fxeEz5mNR9NZnmfz/hQhY7nbW/Oe
JeJCb6VtTPUgeqppxg+zGh+EvYIVlT4kRB0+c0HIT6KREHSlSBdWV8VWtOYw9OL9c0ISTkxCMrep
anRAYba/rwdsUeccaHDVnoTO0rznpeKJI1teUhNC7aHp5VgVeYSLK3GabMngjaD0IhQJE8FAbtfk
vUm7r/S6N20sT2+/P+Gjo4XWtEdIlWRptHivirIwD/UnFflLYqCoWdvWLWAVyml2+/5sCtp7+aaS
+lUsiiT86UbbphBCEfXzF6XrtgsBoldn8DhSb0XNjlRT+ZDHw2wAbzod4Y5nXlwA9roCjydGh2oH
mbmzsPtN2BXOzoiJBxVlWrB0/S/Ts6S7Shc1n9f+jJPcuZGlvsZfSq3AyVxbPvkUZbS0ZoK7+ZnB
UY6jHTCiVt02M0u/2L5Rvj1CXFz+75hzfamgQZiyGH90cBLJHihwj36FJL7o9Fl1qNHWaJ3FBmL9
7rLxplNbpxiWmqSxzGsco0mk3WyRN48Yo7Ybe/wEvx9OurH8APuFER481iyNiXpkmDlYOkgCwlA3
mPvDAdHibPJo0IcCW8nqFns9DzTbP8kn6glr2TVJs1WVPSyRDMek3J2ZB358GCi6CTXDaTTdLNXm
mar22yqjfKg3spaNTj0sGdngbLej4D6ogVCi9wzAvX6sDEcjce+nFmWyH9jwodtOdMm4/iu+8qF3
+6AzdoskllObEYn6zcS5FNTPOvCHpfusCsd3hNzmOt4oLIIG5qAiYClHdZr2aYwnyBL3+OzcMrip
G6jJLkTACnzjvzeX/3xIIypMlA2pBU9k8+EypEY5lmxGzQweF2c4fMnGo0fMUMa+Ud7/oxhrP9e8
b3OfyHETH+Avyd8AEeFYS++zOk7vXRPQiR7fHlvblEe0G3f1vEsd5RoAOnKPH2BGchxPMiqu+ex7
w8PTU5NNvlukRoNeX89nXh8H1XlyONXW6BN8khCltBfOtcG4O6q4HbEb6q3uuz/GJkWWtZHc8ndX
IW8mR/ONyHGLQ8plT01Awgju6FelWl6RC5skguS2Wb7oX4WiPYIjx/JYk2RSZILJevwQz2dDrHcc
l5SOb9BOFohkLjgU4ZQ1GL4NnSNg6xXNWmUOitSEFCYE5MR46mJoA2sGG3k+/4tdX69tsDiET1F3
wcUa+mJLmDFYbslV+PPdr+f4thS/84cSI/tqbRC4I7p8cwQwN6hefhoAaj1cXZQjackJxyuIlDxp
edcgXJutxdvYfUvWH76JTCxfducqGfRVqnRba6fpUWAuprkKVm9I3Z8SwZbMnwiCh2MhzsYBP69o
IRubL420EeTXNIiwg6AP0B5QY3hzYjNXT3GSGllYYt2pfm33cZrgjINNLWgvwQ5cLWd3axSc2OiO
9b47M9MwDtOtZuDToOYVbCFqaNXrHy8642/OwTi+jtFnXo/BewPKMEUiLHW7WG1GdfEXWVstgJXM
ZnQYbPIa5lSnBALYuQ/YZ/LJXZMb9OewZx5SELWTKcPwGGmgKDVpT2LwLAz2MHu5ZCEdLrjlzT5H
TaetXMQFbbdvVyjxWXL7+7LJZ3glc1cihYyCekCbM2exyTkgL+GMeJ5hkel7q4nwvbB7PMaHHBDy
jycq3qkOnOXFAiPy9iIOSphfEIaSedKwOV6aNdiUZ5b/MKV2uQOwPKWhUkmaBBnfFOAEoG96aUJZ
uRFZvtXgYL/o3TJwVRUJbncUWtDV/gnOKZ3Xk8dkIA1ISfZX1CHVgRI8kcFqD3lpYY1iabHZOVlG
3rHFJn6IMqM7QMmjWcDTFhFE4aIbqflPObcFBIfAwkfHDSqhblgNXXETV4H91Lw5FUKnU2ct49Ql
jRMTq3Q4us7yzP4UG4B6LLTOcKAdUWKa9baDupWgww6XwWDPhL7lYtLKU1wd2nREd1/rWvrgwVpj
vSx24DOEFp5JIkTzqeKLe7bWVVo+GuUoagmLdfOJIewBTHx1IeniwqrwGgYDsOEYQ82dbS6g0jsn
/Xu8AkbumQvEPG2a+abIcLRvfYypdJ6kPptfYBvgFbPqYuHe6E/+mzmVYcx+emCbHF0FYlGJuwQm
Z/JkHxz6CcT2EveaN+2OS4G0LwTKqNolo9PlPpQ4PHtWPMpvX6M1i+4FqXvU87w17bwrOyDZ9/gp
Be65Y9Mn4TYn49NiyLMY1TFnQ4Um6IZZEF96LFCvbBFtuFGqOE7nJs52V+OaC/o+nAsKpPhQOg2/
jgm3qgLII9w3IK2ck5hM24BhlhLA+xkIcP5hcoO/SK1ajLAGl9pJquf51Vj5H7Nsf49LDSdznXMe
36ibu0am7jPEJg9Ozswcch/9YPkIx8Z1SCzThHFAYjMNfPMUz/tlSbxJ3E3ZruZDracIYL8oaYMl
d54uC3IKxsR6WWORpfd+6k4XSkFgknAMv1pMWV/Sj9y8jNDZLqm4TiQ9Si8RutIh2C3LPdOHhJZh
D3tBKrV4bH9/xI8qyiaxwFdmwoSS11uUdwtbe/iNY/rpt4UrU2WWNkBYZ7bkta0UqRbmLHrKT+Dp
njtDq6bSUFmjYW8rSN2JYaSK/gQuW3imwBJT36VUyPqRHcjFBqkH+i55uJwGAhotorKWZeaKdT33
GtDbpoF4UdxQw+Y0liDf3cyDxAIpTwq7DGKEUwgTQYAqSi166ndFrkbd5VrTxB8u6h4ZrZzJ4yXp
vcam2F1apVGqFC3X5UC2zY+Ip590iMq5Lgigkp2+71CHkbcnXLB0kSYM6tMTJQKsoueHvfANe4HU
arhR6vGRDXk2+TPEIXIdQCuSRlb2yWcYdfvBoVK/5utglQas0ZX7AoFzXlwpftoHEn7GyxwVxGob
aedheoTKL0V4DXUlkSPKxJbYIzS8BWqqTVeN8aCGafKsfFzT1Mpf5im16w+KGSttK1UpGCzmJEkK
Wpfe4SIu1o2Nn4pcyG4836BuYakyxeoyfMyWqkIkfOIQtaEciH4LUmSIjhFqn3f03OQxW8/hyBcL
tU+Q/olvdaDfG0Nql1urjvFOm2m63EIFOVjuRhnIT+VfDgTfIpNi6a17Rixw4JmPyu04CJNhXwtC
GPPk7gTsopf6r2h5zLrzxwH30bexLxoIc72AW96B6ln0HQPxq2YlnqSlG3xd+JaKM9AhqVw2WAn3
xDgibrfDCVS6bXajncdC7CgrV8T2CxYdgl4aaQ9Df4sVdb2OyyYXt8jIyqal68OhQxbVXc69DN1g
vx+LfPoA7BT0vjg0WIwV6vgMuulfGYpqQeTu9v98nq3Vx+0Pp8ONN5JJgtHOrabunmtqRif7P5Sw
wp+KEsLrYPyuOuT5CEA8Jax7CWgB/BJDYXhE7dtGYxTE+bmLYak8ElGyFGsf8hXhLL1jct1D6s28
0hU2TJ8YAXXZJbQjG/CbS3eCtOUacARj6mzjhe6/hxou5szFHAQzaYWcTqS/lxjHrGKQjOCbjl7e
UHXAQReOpP6KmXflMnJUxvMDcGTsehDXodlgV9Qv0zg4R/TwWLo48tcPrY1ah3594uwlvoN3ULDd
MBnJfM5s1g0ZYLWEZp0sIV/a84lBXG1gMQsONan2jEYLqOyrhfCH68R357AUo0CKp4DKey5pXsfZ
FeuNL1erqEuzXiA2XcQ1DR++Ah83eldlt1BX/5MDuzfWkj0C3uaS1G1mXKZQ5vd2kogXjyPrLel5
I6y/LPlHyAUhqxhaSoyO381avj/kOL4VV7DClKCaTjcUDOXXJPxBzXsDGNA2NnPmqsaRFaQRbBj3
3beZ1u6UsHCcXCp2pl3pj0Ocxm20XZ9GGzk6K/lUZfI7Dee/2/sMvD/T86kzJL1a44rKnf0jX10D
HJRZJidpegIixhLusuquHSB5D299zwNqAnD/AYJSGi91QJGkbDG2STVZpB089lVQ5BbYIz0gL6fK
Ml7zYCPAAVufsZZ75Af+0jQ6zCitohwhl8bBmqIKCuozha0bVNRBVk7IEAC/yuIppV9yDK7cuZTt
nKMmsWVM/vBEpvGIGsghpW/PIRop6hcA9Q1qSMYfOIAtdyGG0dyy0mKBug4hayCsWSE3azHqP7Hj
QCVKB6pgr8Rqz1eiZpnlPLYN1mSNaCBTU+cF+wuGofznr5IZppI1ZqpCN8HhczIbkDCqxWUa9byY
NP4s8lQqgLMUhr9Oq5NIFsMZ/iQpbf4e7wqvhRp8WXLOFvUbkgUQAXtWFnOcfS7O0Q4O4fY6gL2m
lRrMFyx+46LhJ7PgpztVrcg0+1VA3hzolf2rhrb1NQMkKbQA+SU7wUQlx0KUO+XVhyPQLUpmeIQH
NFzo2++yEhcZzmA5KN3U0uvHhrBJkzaSXQ3e+FKY4TKtywsEgQoLIjCiUpIYZ1UCqFcgAna5Mm8u
YdBhxiM8M5TWrB3i8irvg+039/FKfWsBm1BYXhY8qi+qhhvtRwXRP9khabedN23WtrgP5R4wDn58
b3KqFgwsf9OkAAt1uyaTTSGnm1ZiRwAgfyqqPvjzXauL8IooNdGttaeAH+V80SV6ziv3UwwhXAOp
x7P1gGfzJTIGg/uEYFFAFlGCJqUGyb1npQSf+J/cFEaLOwwEE/smrvDny9YllKgF/3ZiSCfNvo1J
PwPzx3GrE3UYzBLJrJbTBmpB5KumH6+oUnTVgRDRM6mTw6KRhqZxwvZI+ZKYPJKviOXDwo2mPpsW
PpFm6ptZi8GO/L/OP2pXnje59yqHb6Ims7Oj2SbufnYpZ01ulOqfB2+/HEyRbd/rMJWQIxZK8sOv
08leaEgiZU1TSNO3X4YhqB8/NZeQYk1yna9x+8gb+T5dHl/VcwqlQhWvD60oOBnvXzKi9WF3iTRD
TseVR0FsAcEEYSiNwTWRTtgtV8NywTfDgnJqB7P/1z5iZaJPMhpJvC6ifnGP1SEUOkytR/Cr3/Wf
5tYeBWpQi+zoX2lqBLMiJfBU3WsBt+ZEzl97WKEwDhEA/KdVoVCRlMwtS4HSaQZpdLTyKPMZ01Zn
x1Cm2HAPbyajP9tIgDPWjTeM36rqHP7hW7JvuaTl7gv1qpq6L9QxvBRZbYIXCyZz/G9uSMrz4yB7
aHsXR7xUpfORq3jRQLgKp9NI/WlPiALe518XVb9nS4RhKsgD0/aebFGfNE7AlZgE0yTAYDfUzW9M
AGDcsqR4psafxyc8b6e1s7FgLAepsvDZ2pox3HuSqOEGj+xoU7MhEGwRjXJ3W3zzKd2K1Iqnj2zy
Xk0qyz5reuVv1UWy/xRZkvIEzAQj47/NYCZQ2NZQwelj5REaA8oAAjeoCQ8VubMqFuEMRDVOfqgc
bGg43CT51Ga70rTccOOxiJrlTUJYRuOS7GkW3EmDOUKYwvspfXTKn8G3DrYaCRG4je+LyLRNKqAu
/aw7tl5C6vRJSo2scWsIxSpZFxy4FmKadk5Sm/IlNTretQ3ogLSwwRDByFryygHzRZAgPiamW0d3
4L3IStEWgQ+C0O4+5FxT3LhSoLuR22UvPYHkoU9JkqZfKquWJvBcDsM5552d12U0BaQRM0wJRt5q
SJQGLOKQc9A/+LeHacn6DPCSCfSlzhnPWB6nqoisW/R+uagB5yaRt0LnW1VAdJw76QUHpt+2HaZ8
pa96IteNa7HPWTOaqAYB+Mll/PfSXTl6Zqq37mZ1d4AryeADZcyaPJxPjnWViMc7PanPU5z8JC0g
sU2s4j4s3Ah7fH7XpwkPKUE/ZvwKJAFW9CNKhMC/UdAnFEn1BnMLEX+EWA8MB6h6HbIxIwexjx8W
Y3yEpQ5zKrSNi+iV7v/zGT6CUUAB8D411BSlAoVnNvWiAA+p3GGDdr+1WUyzb9Dvi2fuMrr+lKxl
Z1egMZWlUdToTyBm2iYqj84NTqpG7JQ5bOnrnLE7mm7OABvdr3DNPbadajyTmFN4wHjuchvsemIP
eHoGSiCvbFrjRsteeOravgvqEpCa5/M3hiOOJpL7fhS9rq8pXQkLG7s8XRa9ynebS2blDpti9HCI
ki2VoJA2NrGs3fbFI13gJL0UH8dyzc7fV7qCqG8sip3SZzqjG5voVtBTz+LSakRGRFDOQwkQGUPR
iZlCrp6GL6cEOmjuhcUCfiyy9OvbsyQtXcJAJ8xIc5K4pSnRzTN9pNe/88eG5OC0z/xivywEwMYX
Kjxmy9mo2R3USSi9zpzGX5N8w2bu6F3lL+NDal7uT5ACnkp7hPfQUn7fNsIjOtQ/SZWZyU9diLJF
+kYOIzrFANsOcw5OcNFFAI351YeAexG4aZjd3dCOwlwQpZt9r5Lh0v5O8B7J44O20ILyaN+yHeB4
WK85P0z/MGjbKRekifxmVN9+eX5p4skAmKj2Tzn4bo7qPVuY229+70UcPOBF5/bOa+aCOnnH3jfI
roTn49JwdhchFet6RhGP00aoLS8EvsHMhE3teCe0HwREO2L+ZNGCEQQnHtjbx5aOHYp4TyiGr90f
tNuARXasRJdoW4Kp+fTVNQxfWCf5hvY5T8z8mWeiHkg6yM2TdmqZhnlBewQnfbZZwynYpNa72Rhg
iZaSJ3H0bl46oBVVrdp/hS5NYpCPWjIHYnxdPje5XAho1j+gwMByyYLUEiZFeBEqk33WlSREDfup
p3VSchQCpBsLgZP9kNmNfrxuwotwA8VL/iPdoQUhnuPCY1fAcZF0AcZeoqb/318A/tTfjvKrr8AM
J3jmmeDel6Y41YlpTPHIkNjDWNoJmZslojG09MjOHu21XQnX2y8ITB2e/mrCoUXK9w9NnAly5xx6
NwbZpXLmgKmnoCTLaXdE3xBlfO3YZvhapKzjXzsKjMqx2udpe1ZC1BaUL6zabMq4ZdUGJzjDvg4O
7mM7IVZGf6RwwIiKaN2FXdNt0BrrW+4g5S+pGN+qgnNk1qL2J+QeEHwaXZFbM41H2BC6YlPE7VPp
3xx9jDBDpPRKcUXbfVAwmwbrgT388z59bzTwmjhz8JwKtFjB5FisS+uR2YoIF0dNRW9V5vCrl4+n
R2HNg31TyknioymsvojWTmOsG0KV8rUTFw0aC+jxW37Z1L2BL62k8Cp2QrT1+0XDrCt4XrrbbPO+
+N+daGyK0ggIM2LO+pftF7OTO+ZnTe2ZlXrUTBtjYgunhgMtOM/O/r8x3e/tPxSrze3AosD06Pz9
2mKAOshVpIOvDKMLvpvQw3vwKB5Za0b0rUHCt/hehimhiBz/4hTHyjA6gcCZUm2qftKgRM7+z95R
x0jnNjCYoR8gobdKMTwEfj2m3B/jDWidY9uWrJlOvALKlAYlRcnZA7VdaSNBy3JamNa19c1DGER5
ROCiQ3w0Y2SJTEtBoEPr3TrQXb6owjBEBvxYETWqeWXN9zJYwFljzT6Hw8MEo5Wvfw2Kg0Ha5lxp
ZWZyFHS3khIUp3mkmTv2IRbyx1TYYgZAP+4BXcjbQFKFVy7PkkGfUl8nRkcAm6PqtVmoj8cBXXFS
WaJP6Ywci69wEpt9vtVP344CMXRVaUqBD6PHJiYwsos7etXJcAynyjWQBROA7OXn7aK1PB9pSaTd
1V9qpx5obU+66o7RhT8xjE582LOZAJVUV4T9JfHuNHZyd2PdJtBjYgKFYrAF8ypvXR9A8JWqN8GB
7VOsr+0JclhEaTqSEESGnVKpDypmEnVIb2u1/h8R7izFU1VUUSn077q96y1OdaSXES1ST7d7OSoU
hcDnEiYn0LqgH9+R2MGDe39/ufIX3nOXLqPjvZDwdERDnwi7Iob+Rg1g0/ZBfdPCnTIJgXKCMaqh
VO75XpNtXyC7em0MUgLGkumjNXkH/yY9lnE/YY30puR0xy7+d50f1W9eOHm9Cn7whVVxb+M7Otnq
VVqZNgTD0Ge/Ch9ff9rx4+YnJz5YbpP2yBfKCpYvjHOMhmJOTTcybLV474HSWZwfxT84o4UD+vvV
GzRbguomiB6l28K+Uftf07altpBIdqxlyXnVxxZGl0gGP0DmnVv9oUR+I8WaRtxNToURIWcl5nmw
R6mlhWbYBP5rSO2G519zt4kvc/N3vCp1FvKKzvyAHBej8enUCtPFJmca9Wb+2/UMz0XF/LuvkXru
6nstDtLcZyUaiDnPTYl6GjecYd18qxOU8aPbh4PjJVvoEYK8rQW9GyydrVchRkNo6QZCgABmOuzH
cvmJyFnvEwEGqvnVdd2aWmVaaOhNKND6mKo5SJ8mVOeB3Jv7mP1qLscw5pTn5itI8o8nwo8vB27m
w0cmqwrB0GJmDXzh8858flnyTKeCgs/titNBU7MCiTHc+GNSxGtfHVZ/HigBmCx/m1Ffc4/s59mv
R63wlSMjK9TIj4hMKxAttRPv4UjGsuuoL1BKIsNo/3lgPQ+thK+7D9MdPLzm3lhPMfF+r02YH5z4
reMlcfzBTso+IBWGyCd5ib9/DJRfhieRDG78zajRomwyOI+6xCQWItyZqJ4KmbFwynm3roeiiuz0
WQoQNeRLJtZd3Qo4JjpGfUpzM6oF1Lqz3nL1Fkt4I5cDdEtaH78LOH8I0UL950cfMg84pfofV7/E
j1qbHH+MhT9ZpKl/TJ+mqCrnjOj14qf950APFujij0K5cne67dVEK0WlsU3SBviMhD88ff+W+sEy
zUBML9M1J0XWOUqkBr1n+LHyh+/FIK3DIvCzGqghBiXEfJ98oQl3AvT9d5P2XmJrzrLJVM5IDMWW
EXM34vUG6UXQOvSLlAY1MMWPGKONA3mXSTY0br2/aEmypmLhYZgeu5PblpCvT8MIMKGt0p6Yq32+
+qbrzQWWADoS4TbLTrYq4M0sHpUQnX+GLNQnVOuk4qdePkC0uHVeel0scKvAHaxxxVmRs5jRCYAN
F1raR6QZ9xhx4fG5JKcnAVxCHADlhHI2DvNSdgSHMgrpsu4GeKWBOf5YEv2Jkr1r4RBDO7LPKLjt
SrgvqiTylKnxa/+cmd1zeehIfvz7kDTdPIR/9pfwM9j2U4TB+VxR87MJ0Rub16LrhxYeQElV8OJI
4Lj6tZ0qQnnv2QSKbHUxwblaAiEhhNpfEormzvFY8krQFrXNnj9pdjKImjLjeOM9hYImbGCTwS4o
hGIGbdzB5HSeKB7hu8HUaSbcAuY4GDkDWCFHP4rmBXQjBoWfZ+AAlORTqFPj2SsmD0V2eVZdv6UM
vMdWlhPrmu4Iam1t14v3dZS+NRJVLM0fzQjqDQu2TPCK1PBzntc8D9mDKxlaJvQy2tXNMsUQIsS0
weZwA75dIepFq0gsl6oXT8i55MGDQ8AH33gAp6pBDUCs0YoWLlyd9FGheSZl7NsPTfNVIqbqg0xU
/ggo+00jKJtjejfVanOSUfAo4JQGSj/h6Cnqk9UoIPVeEMHU81a8xAsYutZBobxZ8jP7ZFlgBR+n
/wOQ622gsS6/AWNzjgKfDw5GqKK43SEHS7cj4uQUbxcK32OLpljbp3VEjMLtFahgX1j51fONrysa
b1wpFieHiTFrOFG+6ufF5rOhToXJpSWIC/1GlKmuSlA8Ms6K84rgSG7jjdCCa3RjHz8ykoOrQ4/F
G0kcr0SHeiTTMbnF6wTmYjNh/2QI68O5s7xAeg68dvYhrcXZtfsJNqdLnWt4qig23TZm56SoDctg
KzVh7m/m2vVsdZq/HMBpmC6U/o4FTMs91ID67S2DpP6GzWv0wxY4iHgjz29S7K9BEN7V2zhRWby4
QYXw6y6QzbybwEZQVrzVqtaiY0L6d4LvLbDfJKMl4tEh5gN61Ih0utuaTFAFA/BuNy7+YSE4IMBb
kNiO0vHWQuSm7NYyonStNiEmNCIAWhWg1/ViyTC1lo1noJ7OBXxX7nbMlm837V0w4n8aWOlrCYtI
UJPQD2KqvQuCH0S7Mqf0pAj7uiPL516FV/BzQnExV83cJxyPS4/9XVYf+YexlY31GjTguMpRIYnA
IEgmSXg2mRBav1zCdc1lX33Egv8zINYVv9VRS0CzDFxsRpGoiddhm2pN855jbGjirc1lzI9DrRw0
eh1ZKWXG7Yud6SRc92rgkCmvJLV95VwKn3mXlW7BzpOPXkHdHfBwqFwnvXyb7vpUnigGg2IShPz0
tbTGBwhB0NZcXjhuVENuA+uY9whD0wzVT3Sh7RIpIajudWJENLUg8SrOZyIvcR/T7gwPTEbtguMG
wMGoCedlbtvf8zWVpvvetzJ5K8FgtEDPdyNKeRNflMoCl/8C35JHLR0Z0UUY9uggM97S0r/coKgo
JqOPuC9/BJnyXlmx6UZ/5o6tPEloFXqSwns23NLIcY6MBgwFSDPG3WkW1b0gYz8CIoPG7hXpEx+2
3RgBzKGb5+yazBYhtwaWGZh9D092JrF3TYY54lILXHrCAT/Yzcqy6ZgEKYpaU81WGwPYCUkRWJZL
sfsl8rPRLoRIbCCgcJG48d5UN3iLR3XiE+x0g4UAqM8chSgUKLK6tZ5f3ZkAd0E6jTsWXcG0p6tW
dKuJLTlmT2g58nekMHcyIdv3AynrOx55qyMM70q6Oobu5O2H+73kd5+MuiTy4A7er4DQNbnlnvgI
+PCcKB0waWeLH2NvjtDb9F9li+nADh+1gZFjZBWf1GtBLgPoDYrW9Fid2S54Pza/dy1gOaWS6hFo
hafSRijHMEi6mKmcDVUobWVMQNesCAz3fsZHruUSG4WKUCx2CoLinRz3Wt1IZczmC2Ts1dHpUiJO
4JQUTBq02rkwyqYUtZ4rQ5Fwlb2VrKqOp8cd5/CxJ8HFgR/MG6BQCj/poLDZ5wthwvtC4ydlv3Mo
l3aaGPH8JWuZoX5HZfm7xellOlgW1chgWetEc2+FcOugjY6z5lxp2akktQzpcqp6cMLCt1b9lnQ8
b52r1Qh2Zihv5SHP1rUi8kiVYXoRo/Lt8863TosSX6fbnzsS2icDN0ZHwz/M1+47eCTlKi+AlNCM
9WKS6CLuI2Rnw6wzqTox407ZQVfr7Qu42Rq4ZNsQc/6XD9y0e1hNF2OUJQyy1WXyaEsUf3Q42p/6
sQwylgYCSp1atjXohfAJOnr9+nde1eJIUzjt+FKazQCentgOXIEOMWrfzEOfV5LLfY6h33SYgd7K
QDH84O5eIvQazjeGhfj9TpZsWk1pZEfMA9oliuSQE9EqIrIXW+UoSTUxMOj2voTHQeX5mJAhNGJT
9qFC5/WAWgksnMG6YKJLW2sjDefN7adSczAuRi9SJYKuj5DhrdfTBsQJU3MpDNJqdFwrbITK/rmc
IjDX99Rclv8JI2TvktEiGmSl5Vp35+aMdBv9xAOOgAsQYUJHgBcdnY7kGzNiIcpqQ7KXPB2029nw
HfaPUZuyzgN/5oQ34JVj57re6ljmDIa2F+MHWCuT5qkWKUqRZSDtZ7vdsXpXq+oMe8putcfdYCWt
4NbAP78dLnmsgragfKHdJBYp2U4J6GrmDH4ZsWN+dZI28MvSvUDM7/pzOHcDeYpFtl9NWpgwMfy/
3OmmAu290XbSHrTdB4b4VHkBRXThV+vTaw4mhZbmhx3wGyQ9UCcwjoGBmm8UkfD5zQNbx4kb/vko
Nrde+9NmuNRlz5zyqhjj8Ct6VkQ5wezZ2AFhP8aEulEvL7uL3c/vmDmtsmIDaGk3SPy0gBZgHi6q
Ya6t2eHucyODkzrHxk3apOkZK2edjLiglcRNVgkoavib7ttpTMyQKGHJ7GGOxk7GQGeY/GYvyvmn
/5HX/CZfhjxwtuZv9GMD4jYXlRFHBSUMpynUMdOy0Xa2qP+LY7WccnlwwXWkMe5SVU+SWfWnz3+g
qfH3y2v5aQmYBT7P5yjtWYhNC/l78JkEzHs1B4vXtEwp00NDh7WS6uvd2QoCAQX1qcSvV8I7WzgH
WdXbZYR8cImx25nALyCQcHPKA7eiGSS3V2t6WbvU6CIYdVHikyEcWxsGppKyfGUFC+GSHfp26dfX
nJrS2ZFWpzO77rbV3Mb+5b2L5lCc8brGczYElojF5IRntoIAoIwx0gyYaMM3ZAde3DfAGSDGs4ow
8igufaIj2X8y2OMkD4XXeX6VlsgAVL8+MHxHrAs2TGLkY2tnsaI0534f7+LpTMqnp2rS4vNZnTGu
oQokgwZDrrfI/XbrDvdPBdLTlYNMKvFuxIZyeY563r42GLn+CN4sWKngvZuVPq8mZt9x/e3kHFKz
r2yEvIhytuhMZpjYK/TLc2ro2sybJzrnhnxAC2BLKr5ITcLujM/8VJgXizJakSEf+JZMJswQ8ioE
6NHiicRlsQwzLxVSVbgYCICZiZ9S9qYGl/OWMzgnViSwLLAGcvc7FdmcTxgo5i2tnx2GEQA55M2y
8Im8BI72TeiLf4qKEQsCInJHwDtEm+Ekjr2jNv8xI+Q06S8cZsP2897v7320DZXQM4w7IH2WhSFq
ZZsQoLQ+bSsFtpml+lRNaHm1rtEjr9Y/HEFMfefuVO/ci4F4TAllO4KvT/P7sGc2KLKs9+MctSMM
v5h5FpZMP5w9rJAZ8R8Aa9Pzrlg/AOhjolRq3V4ikg6iXn18xVQD4egr0dyXNOj9fN0bzC4gl4ml
N0mMuFSr3S1DZPpaUei1e1+/wxQ7VyrUtzkpgf7BKl5wALgmE+54tJ1HcNz6zxt0aSSLIVMukp6M
+Aq4s9FISlqj6/pllTAVhO8lsFdqV2nBQ9ECgvhruiyHDxjsoy/FR0H/A8O4jRuoTg07BTbidItO
AEDUALGpiuQDiQkCErcYsuqzXHc1yz3ahqLKYRb7Ykfi7WJdbmc1eiAxKKgrbJSp2a6wHvIhAuLC
TwfJ4hrTd8qNVqR1LOgrlBRKH41uriKDVkq/Obz4R8PdrtIpBoA3znhl3QHAcxYdcpmik0+T9iOO
HjzP1/vMDaT0WMshclqoEOGGhnaAw+ipxOri0GYjZW4oJwX2LnKODLBwcpbmNa8PO1hwfAnQ5ewI
IA1b23EIxDc8dFqOFW4uIQLSysUBWq8c/JDncAHIVuQzq8/VCpY+aJR8ON6t/9goLYDPDZOByBvq
rbYSTDQu7cyQLZQHKBLPLNUOgU9yDGNg74VJeAHAD+PNMFUEufkKVT1I7f4Ajzo/PZ7rQysLJDz2
DI5AhLgNmqPogRIw/arwqPsDXeRRS8sKm1+BcNRutz5cabbKeytJ0WhVm4aPejc8ZiPJZ5oRaNCN
d0xcJQD3puu4AoDYxppqTmmSX4hrDK9OGgDOf/NU6t9CdHCmUbTdsd0adqVHQUDRz5DFNWbRvxJl
L34xf3x1myB6EKy7yM7QVa9iXR+43jOuJdTP2IN+Ln7HakkgqQ9ydi2lSLzPKJ7Te8IP8ljTHRgc
/c570FGh/4HU4oz2yu0vbGARFt3wg0bHCQS4b+tFa2ZYdETB1WNUTOKK0UbsCQ3Esu5qlfzN9x9u
40sC/ezDt4pncBUa5zmj/3+N6XEf5pJENHyuKxWVHMVFJfKXv5A33ODLoDhiDYVpI6sGZRfjNZFY
rd0fPlG4BveB/CBxd11CEETLsV4H+VX65X2Lt1o1PSPQ78miBcuTLqjhJBCEL6FlrMVpSIQxbeXe
FXlK85quM5tKusldSgm10/NOiCLUyv7Zt4Y6jfpOmCxbAjXWi1D5gHL8iBG/pU8A3Q66kioJDeFl
nAIQXSl+rkGxAtbjxPy73AKhyh9Z3ePFrkIO/8WeWorwQxVHTDrDAG+Qz1RC4QFlRWY31FC4r0Zu
OauBboYlBN44qBGVaGJPI0wvsnQ5Cq2AYLpY/ZgADAdaMuYcTjGQ8hSdJxhN7F6hDD058NJlFQCu
m7pGPWbJdDiVD2hQce0OMXz2FUc2CInqElFNj6BeDmCmGbss16mEuM75I+H4Tx1QzkJRcCMzAatC
BMQ7k0+HIV7NCwVhonqTNCj9Nmbo6cdj2IRcBOSmw2dtDBxDSPhsnKuyOE9aq0/i67gzuLnrCP2a
fRjEbzeSei2tXIzQjTBt6G9ZLctnBN5GOFhqUIGZhGRnZyWlsd0kydqemfj9nYpeNe8cHaQ8ZN1S
4RqY0qFfcPp/KZzx2wgzA7NZ/JSw2Nic4BqmxQxDzczIpjWNkDNj9SGygBLrj0DvsDwwKSgN/Zp8
43wb2wUZyF8NubsfVu48/iY95SIoFQQpf6394WJjXSTx/QHQRsp71rSbwBNOGXqKrR6sHFHE8keH
DaWiPdUUHMIw2RcayqSjNFHBnDf4zRw85EP2iBKZ0DgoO7h6yDQsdEasNIevX5tzp6v/s4x8t8nR
U75kpJztr2CRsO7MQCC9lhhCYcI3lQyONkPXz5hEHaKea0Pd0GYhsvXEWoXQhMzGW5aQLHqfj3Fd
QkdISGJ6aOkKzFInSYrisHyh5+V/D4kA2UManUepon4O/gNlmu5mzEoS6MeB1suubr2v/eXEwpCm
wlBYePHS7qvNH1iyF6EaHxMXruyN2nHoOFcxTv4Ozry88zDBhRGu5G4Nc0U2gpzack57uS8mo534
AsX5pi69P2YTAqblj/tk1m+MEalTgbSnsuGHHG68z1/A8VPUjqfOmOPcUh/lOar5/mWtJburqxVR
TDGsPfnnYVshGz13KSS7pWpdQgzZGUHbKZTXKmgmpurMuygVpCsytfzBtadVXwraavwTzjm43UpH
yYU3f6+cHyogXYFn+JgMUTxqIY3QecUZuZFx7t2mZ73Vy40P2SodFn08fibSuXuWMk0FEjaQbDkU
V+cftC41YsAoX4oN0vDh60sLpTx7/vv54/cPb0+4pEIxm7h2W87zHZwtOvDtZC3eNt0HTeX+0e9F
8jnbdZT/E7RTGxeeog2D5UwWW3h3Vi0lqehuoXhesVmu5WcX5zcHFxmbFLNFT64XPV89wlHJlota
zQBnhQIwyfue5+omz3M87aXfvECnX93VHgNzI1oF+uf1s7LYQKeZeJiCJU1fO0lQFBi5/RJHO7Oz
qxoNtwEX+Ps8LDWrMNhRxdPoJsHaVgnFzRiFjsECaihXzyfvKj3ZGo1i6rqWurN2idp/T8sDdI3s
l9c2ifOTyHRp/XzkTd7NSeBJoFmmN6H5g1hIXAGwU6A+MeO7ndzj/zY6rmt6OABuNoP0s9I9kLim
7ym4BOEnCK3TJOMp0LSQu5RXU8MkRBC9OKqFaWjFQkpA9j7CpLjbVBHVVzYBzKmBSd7CMfEKygz5
0RhckZmrRVImWu98GQhE6vN3vWi9kHHBL9CUHQ9vb143gnbc2dQrKvmachs/ob20ibj48tgS3tWd
sdLZcKWuVkJyBkBG5zn9hiyXNG4VSEDmz4S7UD1jM4azuLVB7cS90IUfXD7kskl/oZwCCqBC+DES
QbJK6r+LxgZfYj4PweOSk98MbMClWoUwhTpZq4DzEsCKQxqNY9OYOh1DfsLeGl0Wxa3ETOMZcB1Z
KM/NdtWQeVfgLvMUtGuPCWGJuXHRJS9mRjSnXaIhI5yOUxwVo20yoU/IlK2Xn48Dw4oledgcR3mS
SifSjOVSg2BfiqYsL/H9HH7AmAJHzfdMKadJx73tSQmZ5a6LOW1qWmzlASw3BTxEJq8IF3cvDjs4
M3ZgnPVt93hooE3l0R53J0QADkDUYSLwQGSf0eM6OFVvz1A7P53alzL3rXvPozQrfZiuVcPNR4EZ
6g4o6u/U3EYCgah3ZNeHtXlyJpwmxjRYu24oDqZU3pDY+SK5ww97nA6CYIoAIGqgnyjrE4xsa463
F0/tmlLjryRSMHQRJZe6mvbeCcY6Kckqz/QDihYSTTgEm5w68+diks9wwPuK5/sLyMiDwixAQC2S
TGzPy4fmDMa5S9WOlOnwjEdTnIlAuRY8S2T7u1qHy1Nvo9dWrQiYhEOeCrAdL3m7lRCBD4HoCH7T
ZqznOm+ygBaXwWcSHO9Dc3zbLHfxebeaFsp2Dwd0dn6sB2O0S0MTer0IFsEXzw6Zs2ex66CujMQ5
W7Yg4okvG96ZK9BRiGn9a2JWM2T2ps2cPTKrhTNlXz+9rrexywf8AsaJRSZbJyDSMEFN5w+w5EVX
zkbxYszsv2ukDS6aIHYo1odgqJ/jpgFfpG3DkFkBjSfpaAkAhk7XMRwDr6LygXht2x3iovQ6kiKN
zuLuOd/cSBGm1jj0v5yU6tdtRIhZqCF7pFko+4WCFUeRKQ01X1sugoi9x6dMthB1/JSLc9fK6LSB
VYwk2wI7sWtY/qRRC0DgDj0unF3ipUS+rBoL/K1MRw9rwjKj3Zqf4MPqcs9eI6mM6y//qcdmcAUQ
jc8/AgAy1d9Fy7DXAbzjhR84D41O1tp1MUiPkjAtLhgBkGi87y7Yd1amkUROadLVcXGyS1r28eQq
9OX2ABYubDtgDZX8LsOZ6Pbmb5tznaEwT1kXUQhm/g/B+MhuPlX4YRrfIaznrjdQW8LoX9GvvPSL
UzzFIDUwEqrl+rIjGxqBbMp9ToMR2RRpH5QzngQmdmxX/cgtcn5QjvbMlE9AxM/XRZarhzmqg7xb
GtDYkOGhLxy5k0zJ1Hg6qcNhZ8crkOosUbMSYvguEY9L4i+9IfaDthQtqLg+hQ/VWXMDDQKxxzNH
qjaV5Wfnk7NHajmTv2TBMLlA1npQifazgJzTwkjEM4j0zLnxP822OamUKTjwdk39khCngKkHSN9P
vvh/y1ZSp6EXDmoW6UyX4CsCFdm/z8NzMw0kR8NdyU7jvvBZIeHvoiT+0pmoyiRiJNYAPQCURcaz
ANLR7pjXdnNT3J8abNZnVmnJqIsHqwSDYD1k14EUcqYtwCkNHtx1czvLqxgnq+KeCY+6v2tZsCj9
N7vMF1mZqwCI2Y2z3KSsrgfLwstAZEML3yQTY5bFD7Sxv33pwPq8Ye5d4SHEhHktJ+6sD5R1J617
gOK3asSSyCuOdMgu2kzEO/uThssaJtuZGINBPze0aSyZ0koh/U0b42zU/CcHuM/W5V/Z7jkPBXXz
rlxfsrKqX30KTGrURHn/fR2XLHJR/Cm+rTvKT6+b03fG1vAxbjEb7XQZmRSrikr44CqEiv8lTq2a
30wBY5eF/MwRuXL9sFBfl59pVW2h6icamz2D4rzY0mg9BuiN/5UjkM0b9U8sPFiBb8FFRHevqaC4
8h1ehSU4fkIKAxB8nwjXdRq6PcASY70KfeP6HX+0KHlz1nNttMd3tqDM/dmfefhoVW3u/Duh2VRN
7ZMg3ziINCsM+nBfvv5YOiPP3jSlLbtApbjvv2lbcH81fxnxkONd9dizltzOCl9h0AcCpfTHSne9
GlAJEb6QGcOp7zcxG0loweu0MrrGoIcbLhkJSc38oAvoC4oSEZdX8HRr1XUZ38ac9xeq1RAG1d5Y
iGP0oN9V93P7ovqjy8L23Z1ohGfN2UR7wS3PZcCAU4Ve5s3FRn48+Yo4gcxE5YrOxRlL/hOhNTvD
57wkk70YWJS+UWZ2QiYEL71pObF/A3/wbHiaJobUvqbBzN7bOynHqrECYFxE0PiUnxWNHNkcEMsG
uJ9wR43r/dzeuAin5nZxMvBU7gpJSgn6vo/3TX/XLIFRBvQ+MFwWl+PIWtipP8iPYN/J3KFHv9ic
Bo86wsLzcrCi58mVuEwdLc4jjPVJfzSDxRagsmfXR5f31Z+bM3iS9DpmftALpxAv10sXH/TOuVeM
SOUYVEsaqWWWSC6d8GIXgLQSir0xB+fYSiFPwbvIcT9q5BGY/SoUJfLT+3WTexB1bMbvAZMeEVP5
EHenkIdoV24NXIBxTAln/b+rBZEhCxzLZRWO2iGyo+vBLumrKheOFksfE9M53mfpqKbRDcogTMT7
k51dKvOzVlrzeQoXHGpw4ZziGU6rhNJqz1GwRUEwcuOB8VWO7GHQfy4jHgwbNK7rEFG7X6Uh1GF1
qkR19hc7G6t0chYm8gOF51rQXSoGTzpgv26q8maqdlcMyawKwdPF102mQ4SoBs8CxxQKznp9zJAL
ssmIWQ+1mnJkEC9b01JieMsmFCdL1+AV46z0sQaTrMtt1S8tYtPEy0OxPdNrj1BZvvh4OP55EYUB
UqeqhBFkWR0NcQ/JTtcI2WYBuHbiO4RuKzDJuxY10+n1pBWTNZpNmhopsAB0JUPOTD/bE7dz2GlP
SByfbqXKqTccckmm3BE9cZaJRX5mdKI7s+4EWie6nnvvE8RZC0OuxyTusGQ9I3nV/VEeiZvoOkg0
qVFWkPeYXk4SofZDnb57+La2hX+i8kKW9XVGq2cafr9a7y/TQpQtj/qGgmdxA8b8CTtudf3V8WKZ
xrNRjLv6BEVFzMULyL/9vEcVZyIWlj8NfXVe7/atdsVRZhco88X3jbrPAOUSBkw5EYkGrN9RA5cy
VHYqPYNSL+fNMHYz0JAc0o4Uj5AMDobfY3AYNQHj7HUNjBrZB/QqSvS6qABhfuryIdFqsvfSPNME
9COCzEEtctQMNrdD4LcigKe7kw8x8UOqn2I4DdSpdQtm2IuPpbv8GJDpERTK0O0sq3gfz176irJd
t+z+MwYSW4zBZcktvL802GDh2v/uHLAaR9SytdPsyOA1WqsQRLMscP6FdqSiUT4Tz/COO8896DLY
sbpww0nYG/43DxtTB+K9f66slgOju4Yf+FjwYIjKZNX12n/sgOPfH+NLx9vug0T52sHuje5KUV5D
TCKe4mqsfhYCcvLn2qH5tIatH6Ujp/iUNN0+IjKxuq329hB/XaPaOgIfQpsPz9/QCHIJHCMPdFtM
7bCBFtz/WF8RqKMYsZATCkTbnl5VZaVRni4hjJy/Cj/KwkF7cAsPWGDfffAlCSSUnMDlgpqgzZqw
qjOxkgC8p/O2BaQlzwJ/S0CoNEEoCsDd2ZXZ0x1YxMe2W1gLyBuD+quNXee0M4WWjfopQj90wb7N
VQW9NWmRcXNCHXQdA8JG2bLm4xsQFVfYeEil16eE4hdNuRg2hKGsvimvBTvlJj0o+eU3sfYocz8X
rwdPyS36hqXrajdtxJ+fYNu6I3QnRbK9H/ZGrzon/WUvR77h6t9tHbHprEbZpvZkmUJO8Zwj9MwZ
uFLUK2rDvXP8Z7QjtXgFlzciKd9W1BzpMQPEfkbpU90i97xc89HEzeu8Yg11IAS7PioK43Go5MXG
rM1vNduyjLNmBOmPQF+dJn8UiaooF8mgFGNiX/LF/3asjEDa+RgUFUHv3SMMF6D49tia95ekMFDo
7gsjt5iNJKQZFcjpoNKKqYnvYjuN2Oprmv5TeqbzXOtITQ2KHPDjUYHqMBu1vvbHYBfPetUdvkFg
bEeybvhzCjQI571wJz9eYaxdqJ8HOWvVXSsgLQnc5cA4BCFeZUyPlX8tK/MSIH1tJe+AZGq7QS5I
3dpHtSmAYBCzGJkvOgy/pHMpy1XwTuexZrru0OO4OKiUxbzGrg7hYZTaf1z52a7Ilxit/qPInGHu
/DVyPfju7ovKhrJhj9x/8BnFvTvhQjBcnkBOpsx+XuPfxGIpn4rcvffh5O5b60NmNTBuoHKbVcvL
/9ke9rfHKfyu+sQb5mkQYHCd9MCx2sdStCrK3jz6oBPD+fkawJq9SvnWXc4xXjbEY5wsilTmBg0q
2kR7+Rwl+d826EXA9X28gcBsqz4LmEigiWXsBLTGWukVjqWwkTdo7dmgXHwOHs12vCbL4MdRIp7q
Kz954md7RhTDtAulm8UHuYd31nuVL/9Agfu0tw7UeFjvOIphCrLNDcCSwvJwhQ2FkyFBPVkLmiig
4ADZwSARO1WdCsaWgiIk9s9qsdwlliq6rVSTTA1xsSkF/R+FiQXX9t/dVGWfuxJHT5sQqU/MytEL
OfA3SIPB5M2SfYx94xTDbEjQfD8cJNqwtDFxtqIKnFJ7drwFVcQ86kpZX/heM+fAm2eIMuIhp36j
wg4DxsiU4NkylOoo12y+a66QpVmFB8vKzfHJ8QI8HjNERYEfeD10kZ+EvVFuK+5woLMSVdkXxcfz
Jg27CNBL7GEfeRh6FBciPAKaHbwbAjGtaC+Ag+qRds2dz2Cx4e7rLhSG4L+PFAONm6YsQMDf+u+U
b1Y4g1djcgjVtFIQmmtRasWrnbvJKxaZLvXnf0xMcg4K6coYKYA4RtFuVxThReDEepmLSKCsOdI+
F2pV0quek0Dq/9kmxSyrK5lqGOUpYMItm4/N/axztAbayPONSN++EgDx0N6lx4oFDONXgBSwhEkd
v4ugaUTGtdTWiCuEPWpsoKfm74cHylitQASNGUU7V1Y6wRdx35foUWqX14vcTyhDy6pkfJ9gdyJT
oETZbFYSBnytJYmwLnA+ZkAijWB0q/mtD8hNsJWlR8X/sAaSbXw3FJT8y18q1XzwRkkq4w7dpb8j
uTbZ3XJtShX2KGn95IoayL+FmKVJbLC3NZlDuzLVg6SVJLoPf9eZFQV+Ykk89hbEhzIi3uiyxj5b
8d9uyy3Zi50hE/FW6gNinO4B3kDw4ojYyv2kfybUShwvDoPeRca1M/cmuhBm00ZYt0XcLQ3DQM+i
56veC3TeP9wMhiCNW7vAXntHGTfX3gvgU+IpXm/Cz8Ta5GWsS9RWrLR+wY3pPA3KM+SrIMmSowvW
chcqH8cCU3JDuuKU1vS2CiEdJL5yA7kCegYhDMFexRRd8OdkBBDwS6S3nXhJacbfU4v6yaozctrX
oMf6n0BGbBWuRy0Zzg6Xdownpv4bWtISPMSrVT+oVhF3o/llKkbid2DpqfbIIinHZQaGzmr0JiVW
Y35XwGkPWntj2iDtPbf+bvFHvwrAM3Hat78nS9Z1e5+V9BcxqtBUxXkeuQYwEn5lFQZTorgSgvz+
jrf1VAhBV8d6xGr6DmX5eXw/06YuUrRZNwqy5dcO6TC6Ez8+orL7FmJ04/bWxDqfvgmwk1XbG0Gq
6DVozQj4tLzYkWwUqF8AHsB+zzCVqnurytagdrfSb0OeLw5Dmw2qIfcwhaG0P+vt/bU3aCBtY/L+
KeTa5XR1Vb0ZoxP1i3QTEfuqFPJELoYmHrtP7FBmgeobAYkGKBupECkrrhfiTKbZnkWjwUZ0upHh
rQsd/n3FlHFtpS8UhZLgenN1cuv7aJRd4yCL57bAoXBuiyN01v2Opee7bdhj4aPHBmkKRC51BM6p
ng8yOxYtn/Sm4SVC2FM2dHm40JL9MsYH+bdRZ7j2mGfUD0awvuGF4in2wndC6V/e383Z/KZLUR4L
g18p+IxG0HWkJQ9oBpro2FT30ajHTJkmNVjK1SILdbfK8PImQ3NhmCb7pwwqdSBwD1yYTIpHNupQ
/4gPuYuuYKiVWU9s2OPj2q3cRMiDv6QjIKLzqmO7wSV945yAoD5Hi7T7ZbhoPGedoAsQmADDPTvM
7WPvy18MpNn6MhJqSdtjmJ5XyXe/z0p8ACTXEmFI1ijylhqx375PNjXB4NvManNlBk4tMrt4iCgH
5ZxdyhU/Y2881kX05KRPbfWI0GWXcKa0+wFgqJW/IbWcvNTL69w2uJByhanzCH/omIkKfyLN18QK
CfzoA5u6rDZcvWavDEp451y5GlqMlJSRoZfcEdY+GoWOPXlk3hIwlIMttlmvCkPODGCxMxlyx7oN
ta8S0N02fbN2WEF0cQ76ghZtMPHXjadaf5Hs82oQulv4SGtD9uymyFtw1ATmrkgZ61E2swQFbFfc
e/KfvcQEhdwZdbHcV5F1G9+p3oofM7hZKP1GdItv67FTbv0aq41qb64RCkNU/1KnhewIINDY+daS
9WVnO6t56xk9r04B6FKeA3hN7JucIItN5kRegMZuqP2MdKxinMORQ8NRSVZ2lftz3ZbRrJh0E/0Z
wdt5O0tP7V+hbCt9IT0gO9Z+Ni2niQoUhhfBCufOyf8eplN1XzShLchffKsSDc5KfbPlBWpQkNrq
/tj8sDC/2RRuYHms4O8zcPdBn9lXlPVIdd5ExZb3xgafxTvzOkLkryvRG2QDdxlWXRQYeVSzf7bM
I7QRyR8fl4YC+CSLFADUjhgXMuppOq6xddPBict+kajAjdbAik1nXdbREqSFNIQQLb6rCSmk6tM9
QbPTXjfri0NQs2HqpPYALGrH/KHvkNYPO9TaCsFLpjdYP93GUrr1LjR6m7/SzapOL+dtpoHG/K4D
SycHQKyj6gvx3HoA4/HodIuLEIog2Gq4mYK9nCJapGZCqZkPNjrQWPRWlUvNlqzdmnT3LlGo0kML
uSOW8fATdWGjYKeHi/b6tvwRFoPJ+qx+iuqQEdMnZDajjx92AJYQo50nZGXapycsdKXQZ56YZg17
bBTUD7pL/w9M6aVjlMtbSCqSL4+7W2d+v5GZRjHd0F7Uvo7+Y5bVnzpoPl8fe5B94dK1TfBh871W
bI6rsHmz84m+/dJ+alIPL8k+SoqoCV9i4+8+/SRWFiKqHKwIvYj3YeOBQcdJ9gK4c5ODTOuPvo6v
ekm93SO174lATjlk8EV+ZO8DBWzWtRGaxNN+HBHQMYor86Y6OM0/mMR7uwRtiO1w+l6pj5GbcljV
ttpiSm/Ap5EA85F1iXhfCuJXHcgxKkZOSYifbzWUFVGKRXQ1/6PrmKiDhMITeVUJGi5/xydwpyAA
YzqwQBAhjjTqzRavEO57lxO8NaOrl44NLsjp2olBwq+0wVJXNzKVclzNiHUIxsHTq0Mtn59mW0dD
xbufxI8o2O1lCj9Awy3ncVH1Qa/d0cx8gddPsRSr1+uCVVcuVywdRplGkmoDfWnOJSu5ipxo8d0L
ACQq+HLFlyjG98N0RQjJOr5pTcmV5XlThtjhhRQ3PyV2PRxmOAZgJmrEvH4dHIv0rwHc1K2Dprdh
PEtf8CkRQWrQEytY1/1baPQu8GT4/yoch/gdu53PnJri5dBf1foZfp88uVH49jn6p5pChMlfj+Sq
TKahoCie1vA7pgwhMClVfy2XGaM+oy4eUhGW4OnCEFG3QdDnjCSD/NwN5+9qiMLGMjNHDbdRMJzX
xZshuJJCKI0PZ0/phDT/OHyjJ98aOgml8pNDJvpeW7kCH0/RBfjpZBJduOmiN9mWwhD/MxoAwyrS
5/6jbhowvW5HrWFoTKzvLZ68SdSfL9LtSb9Q4n9hLnKyekRHzFQqcCwuaPU3aP76xCxyi/a/haUx
Fgew3V8QKrMRp9+C8ccpZS72nzU6FwYzz9++adibO0UM0SlUQow+8Hg6dNhdqu9DX4hA6ElPmgWZ
5vtA2++Hz+jeYHegPTDwlHk07nOQTbJg+gg39BuAjHqw3afvR8PXjaAHbh3pD3ytMheyyqEgh2Hb
HMWs4nrfySuSo6cf38+k6ErmUm0aZx76YzLLrb0U4LqeQX05WEMAfMGrUFjhOsngxtqT6BYqFvVb
DAwzcdB8YqsVq9nhuJ1tTpY2vX6jWe/9siMzGVygw3E0qO5+RDwtFotBHeRofV/TCSJlPWW7uE+7
MzYp5+Up51VKBE6lp5p2rN8r1W8yZIVVSdUviSHNe5OZQrZmXp7Jmzo99Qnei+Q8flllkYC3byeA
Yt6GpZUQUVm3pBOcXm++DQVZqZFOqvsTGOr1pI99S5Q6FGPC8MsBQP9uD9XWPeou/nhQOgdVfLtc
87cewLjBqIXSscd/ipSzXizB0lKY7av3QbqtAnQncvXXXCYYC+R67lyYZ7CsifSo1CaVpXIhBoWE
rp9LOzWNMBcgtYbq/uD9BV8eREd7P+kCuedolVez98lbpmog0gyWd6ab2XqQ+UHgTMNfA1HN854a
8WEiktf4mGbLAYn/610Sk6+vs1LWX3InQ1UqPodQQ8YFAu9LgnlQDUJj+ngdB4CQOZ81hBO/XnkS
b03bIJxZWpN17R12nJ4Cg6idCimLLZ+j4LNYbjQl4ftqj4VI1OAet967KXAFtW9Li8YCplZEfNJc
3ts7D7ZVe7/ranAj3H4M7ecL4oTNiRbn8x+w+mFwQzuTsrE1GzpOCadiL0PkPEzlBpCIvxVWjOZ/
vPNmnFT5Ci+92KClU9aLgL9vOcLI7JmDDrpC2+edP9GimnglAiIJHoUuLuPZ4DmvcMiIul4O9nAV
yEVEuxXoXbwd/feG/sR/wlCRqusTo11HWnlBPJZwclUKRclhJJ78/yHr60W3mkM1j69fH/acJqmt
6KM1qAdR209PgMFcyr6aqhjirzLht3H1Tfm1oOjD59Dn+H2t/tshgCQu/aT0oijUpNN2F4kukRIz
g6mnSnPBPXRyA3ZM5NMKKVFtSC3xjgA1wcKP71mwkUaO9rQ+IULOE4Y6hPn/bGkquY7a/5w8ZaNB
UxPOPsKkaT+6GSbsKERWhXO3QFL7UYg5fGPTm3hr9iIooMT4M6DTOfRpgB3qz7OOW4TBMZDhqIn8
ePkhDq0qw8+W5cTcB7RPihYlkClxnDZtQjmJn3v9hw0//hvqAII72jD0N16s+4KanOK9FAok897o
JZJA+AMMI7JgengvonGaiTpuvQqeKvNfojo67KTPPASqO0vZyefPO2aWrWtyiubvfcfJ9Ot3U21K
wHNUo/yJTv5Gyt9qnZ+dAQpBTHXzKQqmgKeXcMOnCDvUzwiBAaEZhBykiNy/b1pxIve0kcjlfXUZ
AVQlWmKN1Dp+OR2U5XIOY5ULObk5hqEbuyXLxlB9VMwpg368+HgfF+wumnomavkEpgKgBkJt6AaR
avK8LVw9hzEQlF6APcVtRuOou6CcUkMLKl+3thF0CWZ0h9X+4JIJDqpxeYEvP6eEScEeT8f6Wv8u
95++c4IUdoXgt0QytuudSHnaUhqblsJMJlzwZ2L+ApY/3WIPb8lSXsOrzWC015VnlccSvyTOm02r
BthB6jG1m+MjXNQ+Dm8Vnvu3vbftAssQ4oiN0nAkYE41faD1GiN9dVOUBxM7IvpSNxeLUuwHOlrA
b7zekjWl9me0xtsM97i3tYjo8Un5KoB8xtjjmMnTY/pMgZZF9QNqg6fJ1quwbVbC+3zyqUZjMkt3
cHNuL9lG4y4Ot3lc+QGIOy2sWKQl8n3uURQO8L19VqYsXdmhuQJiyZFixW4LVVq81rQF6A5C6LDx
rKAS2u8tgdf7IoH0Uo/Crb+VOZNtQd7bJhmAwXGazcltkHELkY4tPwMLJrssoXUHNVEKLmszKgdh
QPb83QrSgOOtGP+NKg4HFvAohS4msOwVDXGIzTinvgVKKInX+n1dXJwZWgovlgaQrrKJrxUGPoZk
+vGgKeNU8ZfnvRrciUwQSEAi7rYAjakusaSsFuV4Zh/Qd+Rct1SNtfoyTWxNbtU8l0EiBA/FJXNB
lRkBy7yGiSIQz3ESJH0+nxrQHNxbuN8Rbrh6yc/aTQIUaJQlGfppllpv1N2QK5Rf+4jgiHYh1l83
5ryNa1FvoU4rmxeFYEPDsf5OnKCZCvO3SXqPDV7ky1VSBh+bwva4v2Y1ATDwSDi20Y0N6DuzGUZT
r1RhexY3qi5miAzBgTAx0NRoZpOpbXIXR0UF28oGL0ikTNYEemOFe8AgQDCVnkdx2qstMJbqNheE
ZurktgLM0SFgE79h7eTIYp1Cy0qu0gvJgXF4x0GEsecpWKUTwkT/dWm3I16jsA0ATa8jPrm08QGE
2hg7qSnzHLIro9YeuIyB+YAiM+Ig50v71FK6Di9GyBtoUXmETkfZj8n7v/M+1C9wDq5eTE96UrEt
lNpfWckh/n9CBJS3vxuTxux8WYrO5AFFTfolnfG48aOxymWq08bc6R8zbgwg0iARTCHPijZkJKXz
pK/ti4SvQ3mkVoAbQAGkdDokFHVdTwepqBFNWYoZTINt7RGGGtPy/gDNewc4rqjMZrQL4ZsFgCpt
/Io/bJo2i8CzGd+/YPqibTRjRrsG8q/U2fOnpt3dU6sD+HTr9KMW0z8Ku0z/A4yFqmMPDVoD+Om4
AsgbvsYGnLGXYyLCkUvnoO23l3wQ8RJ4hVBhf1Tx7hsbsTVs26X1yc3sKWhXC02VJBS/aRMTrR30
GZ3tJUCcK6qva5HyjT5M9Xzw+dSFN0HMpBk2hxBJuU8Lw+54Fbuv7sLR3lM4EJh9yxMhGFZ560vq
WE3qLMJxH0Dqj53xxfTTiCAs2zhjkDsVzNvkJeN6YQxfnGewmZCt4VPfiCsYDn9+egbgCxX8qrRd
9FP7mtOiUkYU8jvffgJQ3Wpu9Kc+vN4Fw75bW/LFALuyS5WVDyih6120TE9yZMYlbgyZodsO0+A1
V/E0gL3L3uSmpQaHpXnm2hJjNRmjoibkzdSiYSaRaV8cgCJKUd+XucLNo63qmhEhTa7xy8IOrk+O
fMEaAoNf3I4VGFrCujWfLUevwUfIGgbJ8REh/kcSJRHffRe4/LHVUaKGVF1qM2IsSF5ENNqjWU81
+j+JiVkpLUiqJXaq+j8dAHQzG6xxzxt6vag3SgRwVgbnwb/vO3Gq+y1IW+QCpEtAJgUV+GDdFZDU
oObQR69lKR4x8QtN/mU/QrXYo+yOno4a7Ky2K4nWa3svosf9e/90cqHx5OpFNtivEZjM65QJwWBa
9fkuWbq+9AqV3S0vJu+3E64zodmwKYLcY9mxNCiXx5Nn/yyNpXs/s6xyvHXGyvhMbKv7UpgS2ruy
2CexOSvvUZfIGarZGgr8ZTPltGb6Fzj36wabBArV6VMi7qmkmXgI4Td+urLgWjPx6/KobDTgHWUv
nDYnmt6T4AJoiODIftadxwi8AJ7Xl/rOkd6tfGTDb0yKbUWyuR/oqniddOWWcl00ycp09XSuRPtt
pSY7qhOGeK+hfJUMs5xdjeOVblfS7InP5fH/fOSM0dNL0Ksmam/Y/s7+dlQOO+T6QUGRcaqENUMk
cadU0k6IYPsgzfBN5+ri0Uej3NPKBDD0MZn9gT10ddE7U63sOKXgAUI5mVk0wjldPmeXq2eTocgJ
VLo23y3zgx6LJAC3DdRXQXouVmzsHwWpoado3YwTkRwedAazkGIytj1kqxZb9FMFXVCPXbvLcM5O
+zcET3wCRIj3mJflBFEg9bXfTvq9lNg+sbAozOUqJqMCoQjDPx4U0WdCsw+cgfDsH2wTGSSJIdJJ
n7QwxOMmEX/sb65CF6lvhJf6wtjt3z7dvwu428bFRv7+WVR/nQBoPvKRPD9+1px5aN4/n+PT7tLo
aXq+xnuVYB7E10Q9Bpv058HJlzzI4foG8DNGB1njX6FUJ1V3HnZVmslrcZxmtOb78kOTx01EGlhk
f9Gzz+UM0xwoCuqGdgmK1mRk6AwOL/xbQrdIDbKavsj2T8+TMpWhkFhieyox8YXePURg78jWmYIM
EvxSK0918068e0SgGTddqvkTq0AHPMSkRHQOV+9xeQTPayyVcZdWGm+iVSZmMWbZV6kBQzSv5cQR
z/5rIARsf+rCVjjJe3eFj23tftFUqm54RpB7X77Bz3dRS92zbKT1gVOVnZwTcXU26WLTn+yePsAy
F22OWw4xZJ0wuNkk+kqMjooRFsJm9kCxSehJZ+VZtBOLBnXTZN5bH/CpIoRp6ivRGA3m+b2z8lza
qnyJgBpFoF4a9YYzB3L5Xdw7DxHT8P5EeZsaawEirdWfIb8+wxyGQTmJfcUeFkS5Kp7IO39M6vec
WGXF/5lJ2//sG8ncrGvpP1KHDHLJJOf2pcTt29UeC2od390fVSyC6r4DAPai9jKEbLA+Pw0Zj6TB
DrcLQQSb7tbqHoq3IUD48QuarRTLSKhspMqb264QwLc4MoFvMYlUgjEEuPoaBWUcKMyU1UW1KVGm
JKgvutc4FVE+pu9EXAE8STiZewr/LYCIRjrLeeOMccwsMMgIStipp4GcI5fxrS8Vch5582uLkrJu
JE6Sy8OoVHp3BaNnb4RPr25AfDunJeV0+7P1dkpr06VPyIhcOXFZpb/Lsi6JQ7ocVJh1fdFmFrHd
PPQsxKBTycHBHxGbl7qrM6FANxcjqcHy+NtAUkbxG1FTxmberQAqdPDhEU/yg8abTkGAxg2oSwc9
z1YBqac5tOTmIRElnJTqDCgm7OXfHTR37deyjPVdYtGChKNhsvCqpib4fUoNCPI0s7Ko61GGQFZ0
UYdei37I7ONelAJYsiwolCwLoFxRAllQOp2I+PjwgOucDQBNWj321oJX33ESocWAOnz4u7RCk05M
up2xTTMSBywPaPwjkkIzdcr8Yz9/lCXMPUPbGhQ6zbaF8lB5m7IPY+NOMZAQC5+k7HHd99kXBARm
VqbJvEcgV+CDABs4F0aKRoEJ5wvixM08TnHo5jXMcJbPEgSpNmc+8iBF4sLzrNYKKQeR8hFpXNOM
vC/D/myH9oBm/2MwQoDhwF6VJI910pJyQQgraBqlPB7jXSiVx+oqI2v60Jz2jop0ERc6DhYD+5hc
EnYINpHQTEpzYMJv5xlUKwIL4U4qpliNaq8hijwPaIVh9xHZollYIn+LhE3nOPauT+DQNMbfQBKy
oL5W1GKI1sgtIA9nZRXIaH5Q7i5x93TnkXKRVPxBSAQ78RNgusJTIdvqArbJ2/vmZ6G3TLC8FH8A
Z/HFlogim11WimVNHOTgAx+eJKBgqvtqwLa/zP/EMHPsN+Y8UWXutrsYuicNsyLFFET9hNPuCROC
7wE8OIa3KTi+EEG36fj2AioXTl3jDR7wDBIEfZbXeMiR2pIjifkiId7MLlCnSY8e1pdak8qDAVd/
v+SasIiT6ZWK+lT5WDoqtJxJEGSnxskV27imcHcS6+f+o7qG91GRX1h0ZP68atUdTb2YIeNZ7OlR
Hq6ynvv2zFYGSJ0MYALIBMOviinoEmICusZhEYQNjAgl+fVuBT+PWm6xNM7HWXpeQw6uZTvU1g7S
rQjyTjxHzV4S/a7WqEwVeYs/6DQYQzLFTM1xaoYcCbTcUAWwtKXNN2FqgV7zda5q826aDXeBLMyW
je2msHVfjQp6Fh9xUGXWV1C3e6fYbUp6pHiclvPspIdzkEiBVCDL7LoN3+Qt/TG/A4ahA5rAUtEM
Vj138ge1b2WqQIfNruMi/3A5v3CaivWvFAuaPAd7LMApBAArYnt91qA/1OoYZD3qQ6sdpPHlSK68
rygqbvSeDCCsfcAXtygbKO/GpjjsRVVFrjlWw6oEaIha8kJ1kOL4VRQtNwAFJn+ECamSLlwMsnGH
Q3+flg8AZBs6BiEsVrqaOoJEcoDL2aGZOQ69j68J2QQjpK9D7Iy3gFDyBhE+WeTuEB1z94ArhEYx
ParoibI6uolA72jvt+POONUuEAvCkviBrzjmP4hkzFT2r55NZWWnWkVG+01qYAvzR/i7QH4wdHaO
oy7CAy5TC3bkgMIQKizMSJoCqe11tMhDtiBYYV+MnTYuYbl5bXraIVZ2J22KRuP0a/NVfEHxww1w
fieLWq17t62PpI1S/U+EPw3xOc8Zds3qxjor/RB4c9OdzTJQ7DrhuGlFC6ctbObQR+FaNOmCyt8u
KPXqZS2abPyarLTDrq2Zj4AQBhk8tWnskACOOpo2E/8OQKNRCwyYvahn1ZwpTCMHh15ECHVB7oKm
5QPFv4JfxGf+u57kO7DBP64exn65w7EZPKDM9Qpi8SewRkyzXP0lzsowuikrKh9THxEHO1T84Btv
82KatzVeqwzcozcDGqcZ0ROVBQ6JgTSoe6UwXqU5tsbDURJpMzD2JJGkCwVz2mCxZpD4pexp/gmo
2pQWSHuhU1usaiofMGMXAyXEUbN1A4NgHoLWTDB+QdPNw3qgx/4Yme99AKbES05kumGVsbI5vZzS
AOctAjbUy5ur3ijPdye8ISBuUUaVCIJZyQHDjmauxdFFDJ6huX47hlLCDgouRyieminj4L09bjXI
8/gNlVa8XkMp6j2dB6KH88wTurPOwozYeXsh12DOU0j4TWltS9lxtQ5eU9luZ4Np/cmx7J++QKKG
g6/rbGW8dFHRWtTckPIbfbsG3a0anGM4OmLuCReVZ6qZEaBcgfv1lVko2KzVfC7KB6XaLiFd7wr+
X7nnYs5O6elf2v/RjJgh2GJw69kfzkoJ8h/PZW80s8u8r6kHBttzQvOXTwczAkYoP0r1GF+hrBtV
k2l6U2q3yAs30SZPlkehLhByDxb1xkU9ArBUs0UtuBWzUz+Qzk9FojoqlCM8NRJOtqEcuCxaRM+C
5BrPanf2tq8m4EglvgiDookWKpaeOVtsZTFLOB1Ui1rtfjZJREuBi8henF31nGRpLOQFZzRJCh/+
JhKb3zofrR49SwdvlNfYdurIHIcjwhUBBiJP+FKqCPvdzV8Yy5G2MvgU6Kbq+VxQFIuDaHyI1feM
bt9dZKdIKrVskPmoCvMVtO38QTbO4PozXiZVywTY5BM0+XFUEAE2QPNPpW1RUjQYlPu2Bm40l9lE
hBDRcEVFtH8GqYdWhUZQoq/pNevhMZvKb+3qjb9NNCIYNRrc6rZi9jfT3ctNezhyF5wBZ7EC1v+U
CCDlPEjigczeJAjkx71PYLD7BsuIuBhqWkN2UvYb3KM0j7xNY3DPKBDYwRxU4WBhgqMVztTg3o5v
2r21R/PvHEUD317U1a2gVBW6jjJaXYLfcBQuQltGB+Emz9G/qc/ccjBkj239frJXKTSHGCgUxYmJ
2Vl06uN4GGcfr8Z22KT7pKP+j4zMUjaXLdjUv9/Ou4O9euEz5A+33xnrnxZDfPvbhTZS8wsZhHRB
+aFRiJ/IZuTGxdVlvg3hqGI52YNKdntt08UcaFhCM889mZoaPvsM79fdzGZsJmujxcJulecLK8iA
M+A1Dv5BxMmHJDJx4ACgMueqwIwfnN8LaiNs1NlcC7U0JurDe9NvTNSn3981uqaOjLKPGS0k6R/5
a4sLpqDd7iHwf3kWW3lqDL9RHF5TwzZuieE6JRO1o1xb1suMLYD1G2zx0AAQQiExONHViTqmj+4V
w8Q5Whb4IcMQAXHeVEfzBj3MNsYFFZKkIcx539XM0yps4YMI8cll0uwIjSzPIZ5ucZaax/ABco/7
WZgLSt9IG09RYfxD/+Ol7cVLgI+nCYqhqth5B25kQwnFwGLT61gqCWv8QU015Qk64qQArLjlg0ft
ZGB2IlCqpEnKhx8C+pCJRzZToUEVtOu2muCHTCJ/fHwqAJ1Z/ozJBq6EHoDz63Ym6p6//bv368SD
4Ifkm3adAFl8Hz7WqOupkSIg3QoBvdpKnhcr8jie2wjpLKoM6lpV15pVcWZf1b5J+05izbUYGQFJ
+RRmX/nthnh258/dQ+QSoaPGigmNHU5AMGuV++Ahe6XsnOsMMTHnELhlv0Gisef0cEJkieoORiFC
Spr9+hOtEUOvep53ot5vbwOgAQ7oHcrqy5YQvvGKOnlj2puLAXktIUjwPv1vikbRKHD6zIg4T1I2
6P2/sA7Ron0hJKMGXe9yXAvipX1+yUU0OZfxem8kKjLVKLdO+OOUH5w0bn9nzYBrxLii9uq3rQAu
fLcZ2CpBQVCZE8s3/2KBnTdRGQnrmUqY9NNoJQCMxWbmlG/cnsBsUKk66W4HmObuLwSR1UaTycju
d43dGfU/ZthhS531g3CLTxNe2SXPwkwj0B/lPjViayesqJTlwGeD2uSXesLkxoFyvr5qoiu/0O3l
FfEQ+fk3XD1Nxe5QRQlno5rY2PyT/5QIlKEhO3jFPK7jLZi3BZR24wgPZAlpa7wNYoYNsnQWyAxO
PDwjGGYgtY2+DvNka8sGfxFeWmsFePoqja6LBWn5v40VvablA3q1LjBCqTbuGRpCA68+BOjZmuc1
t73130ckQT9WqWQbjXFj17XuiJAzbY/K3wawnQLzVBREkEmpoxxBfnHgs6PgnfmCeaMPJ6pcqZkR
y0LVW488+RmzsDf+WeCQM1m5H6fF9xBnVCQmH8knC1rlU4sbMc9VJg5UA4ilPie/1ujGA44uYfxr
xn1g6OaI5ztMlAqVuaMz4Bf633wGvHGUsHRY66pBEtWM69HpluRuxhmWd46qYFs9khl1lIi6eWCP
s2XTM4MwgFQjbQ9mqoKdfvoIw/SQSxEvuLJXT9/53oKGklgS1uMPRsSVva1//XOFmAfMuFdHUsKg
zpfceDDERVGF+kXmUtkN+WhiPj5Idh7CgjJB8edWqwYaK0vkT3p+n/iRB5S8RRyojYRXa3WA7u2N
+bbPACl4oDKyGFaHOnYV6zZK6w0a6KkGx6BrqkwdXxnjauYiHbFB2zVE4sk7XdZYCo4GNn/4hvFn
rSszN0TUJoVr+7LyraifYMd8oZ+zuQ6aOUWCaYO/ca4LsUdxewNn2KiFV3Q5DDXLnl2g2h3pzCzD
ksXddLhHuQ8urpZlyG7+81It0Khp12+HjtsREoWMIq5vFgcdcmmW2rw2QSi0Z1MgyGa7PQ89Y/8A
tI9rDSBzDqip6vCvxZJm2YFmcPoFY7bUr5ysxOJnpyMdGmSlidsBwH57G/kCJjcTiFi5sbihk++j
qx/Batg3bXEoiZLK21GDK7uJulfXIsQ+PLz1ln1t3opMEgtfVZP4KgQkqjOPSzbzfRNNHssqMRPY
pkWiSxhHE9BqLj9q7ewkIlpaPcLrVVkC+IS2I5MU8NGwAvjeKXiaGvcS9RSknzkn89BAwbIAuDoB
0L6PpZ7lPZ+th4n6oMZQF0iYGVEDoD/qrRrzFg+Pi6bKOcNW+jIIHP/q+wTsvtS9Vhd1+wZBQecf
leSAe7ug+KZMMfb7Z0xE2v/sYOsKUxh6BQ85HIMENjVQXbt0iPwx6Glw6Yur4vGeMq4EASpucThg
0ba4qYIAUMSryG7NqQenynOqSERK3sVgqNTieTx6cVXEyc7oQCzBnPEeaJt4G5jo5BKkWATnI7fk
xPIx7fiOvr2w6qLh6bUdjqkXcZ3YWdkoT0cVuIsF9mPpaetXQAkUV/c9W8MALCU5Aiu/vJ6ptSKI
JR9BsVTbY/1kdmbooGrFBC1iWaI7+XDHi8nxZJ6wOgD6mTwjPYcg3dG4Zen3m1da2u99N941HeUw
mkhkhOcMDN5hI8ixUZYL5oRApngfidBAJxcdpvjxE6JA8iIAeB2X2qyPXI2nxaUAsXtTUwphJcUz
poSJgiyAok7ii/adWKGhmNt85XidbYfNAmV3JO9nhK9GUkHnUgMtMEMXa1K5EykHCNeBD2N5pHHX
SBq/CmUB+drsklyyVIlMQc7XI1s1GddHgdsXkg0FbDiDjnRvnMQK/WhvQdSbRAApcvqWqIybb9NY
CgGwl1rh05qh/FmgCL/MTiwki8t6DgGJlJoGKBDc2qLHWv4itPxmy17+AVHxD37hy+JRDPcewYqn
/pZKzS/zvZZ3GcARsbVzyXn3kp3TJVCssUWLNCptoeojjLsfjpWhPx3l7Y7YUXzvQL+ibmDkUgXD
t5hRrp4die18A3h9xQJoDQT/vndwBxUF7dMIuJ925u6uYUQrqVAMwriHW6JKbPm6KBkoPvrdIlX0
LW/jQ/KM5liyTU5u97rcxBnmO5OaKKVmgOZ4kYT54++hnv/CPbBeEMvfcKZmT6pc8LM/jHDr+4Qw
45Iwt4+C1iCQ3YlYSVWdJfVUW5pAB5jvnEjR8K5k9NF2WjDfoDhipXeC1Bh2NSBGQbweQF3NFOz/
QaIUCNREEEaYs4JM1zp4GZOuPo/Qg2vzHx5CpqoIyY24RRYEEFjCgkoKDdf4zW7QXwWlrd19HOBi
4j39lyWSfdMWq0GGV8caSQiF7eHRUdE2YGRxwxxk0CvVyFeT543Sv2saCpbQBgsbBw1exMudvTOA
dqxOynM/Hn4mXChVShFzcXCfM9EEEYLRZGMxq8OG4wgXKvZzNne3FmGfVTJ8AbH8mWG1LtBmaEkT
Xim4eWtlGh0l5AII/0A7XvyjAVuFw1bYgehgxmRzTSB0ztBiKqynIEuFiWiEzxW0UB14E4myEpJh
HxPLMgDZ7ArCljKihnTAqdMw+Hu1sVZJiUpdFNJwaoKMmLu0z9QvPVKUnhfENRRGDQ3tM7duiuzV
hn23IwdxuwTjxZl0zvtFYrZ7sz3UDIUl/Y3LkU2JIOnNFGeKf1HN6tzOXir0CnQYjMFVc+m4U23p
KN6MdEoPQszraAT6Px2wgINt9bzQ1ot8y/T0E4cJMcPbF74qQPi5UsLYquW6JasWoFxVS8GJ6v7q
l/q5rT3LrhAHWjDAGcvoACejq/MBe4hLJ43y3t5wkYK70Wc7MT0yX8bPA8eZHdPquWNdnBG8v6pb
iXaStR4kGg98U8Xeg+nbMCJicPZpMw79XakrKnvSIIIidgBGUVlPVMwL1mGWHwXDoqS/7we8fLJP
wo+5IaAYkfKnfVnN0iRKw+g1I1RYCLPfx66n2jRqi0+dqOhKJJxqX1tNxRL5bACpAfigRT8heTQ+
ECPuI9qPANXHWdX7lxL761X3KPKg7XmbOlBCR8SqdbSNKYoDjgIJlz/ufcF1jSfZ2C03Y44sMGDH
85hpQHsrHU3nlp4XhVSBRS/SNjSrUXV3ZGP4ocD751P7MRnCAD3DULXbZOIxeJZr29nDye22sSjv
4nVdwZs3CEqB80O4XrlwX8qN0nNTWmRP26BNBv6WUFaeOSgUEMmQasQfz+kRCGjYx8Cx88Da0nB1
GJt6R1OxsUizx1kM6gLAjzGNyLEn5dm2pE3HPu0yJHydctq97UK6FMMTNafCifpaspYKs4C4+aTR
OMG5eEImF3AVpY9zpuVhknp6Nd3/Hdk2EHm39T7ozjljOi/M5/JU6S2D1O1tnVuUmXKQV+FyhrLV
GEtTmXRjNK5uBJR8rrxei27j/J+m/TX8FQBREQ4jdnQEz0Jlg+XMVCKX1JPAZGn9/SgfTY/utMxJ
gL+ut1ZwbSl9SieIUsdji6P2X/BJOhcgovSyWj7Vk2UXivMcJAYyrFYVrHxCKqOkW0qcki+gYgHC
RyJ/fMtRP/c8JuAiC+NWlZ9rLDrGAviB1Sc2VNaLD89hobhF1JgqFzl64nTmKIa/FgEWJReLgwGc
+o1/TexHQ391RoHrbCXQAzXnHi4EtpiXCYdT6DF6W2kSYcg186TIYgvQCRkiLIIP38MXBKdiqEqO
emXCjg5SnO3MyDYMNWUusyaIB3Zg2urNku6fLkY0gezPtHXU3htBWGzwYxuBdiotsAyBUW0i7Ird
GYC3UC3BSjOIOP+76bChlgKPiV6K/5EYYsHoSYoo8XwNH24fDVqDhx+cr61nliPcWOm9fVvpB05g
qaqIYvEAlzwmPyxT5li8KZw3Ab5GuiCqKqZdSAmXoPlt6pihl3T5WjtqR1YHKFecpDmRP+u9yUju
WxAvRHAdOoWCQZpa8q30lvkLZkop0MqV2APrWV5s+99uOzm9Yr9dOlgBjwAMwXIWXX2WFNT6oH9D
cPjf/ZkUEfMLaQkm0rruQO69i4lzb+hnGPk9CcnuP0J5OYz8Zgnw7cFcnxOfRxs8WuptOxG2yeEW
A7P6reszfwS8QGvcAhFv/0XVFtfMBNaB33zjUU5rMYGdOyKijojJ2K+Koc0cN3cQOJBFrAGagI37
hxzWXNHqXMgOnzdXN19kBma/uupOaRUNQ4DyPKmVL/aPgrwA5p6N5kyNsuK7NkIR5i9M/QU3CC51
Wi8aEP04P6lWifIWeeiEq9IKcHtrQpU3E7PXe5rrqd5sGHWUjHgF5cVeeQY5bRJT5o3QqJ8seCTi
8/VpqZdAdLr1UHaPUEAgNe6mt4XcWsWF4wi3nfQ6rBMQZQ5KjEQ7i2KKVUDj4T4tPDqUCtE/SYKw
hHNgdLr7ePCx0poae0Q4VDwRg3cGU8cd9P4pRYVn9YQbTxnziHyWJvMqF0mxJzSTjloEsJzWbrm0
V9uEg2IR1CBDnxhEKR+eweXdYcUXhVPw7R6zkHZsyAyiRl4N9BYJXj84eYATmssxUNjEWE4Gubfg
lY/p+22of03+a1zWkAq5/7bTbMPhs3DUjfvPM2tdQG0i4FS92VwFEBN/xlU/qY8vzoMcIZR3+eTx
1fId83ZlkXdKwXDqklJu+1c0nfXD1D0sW9YIxejEcwPZVqsyC3Bkj2SKAIjRLuOEGzX8d9J+ZL/w
i5MvbszpBOhwLKwdTUFiCyY9tb52LjyAN4ZdQoCS2Gs8ZflWCWFWvItsEXUzmkC41kKunqvN6aVg
Ds3maSoX/MsRedgeRdyAhlPFUfL4RgnLCePcV3uZckhmzFB3tFp59wxRjIDsbsF/EoDuFruebqkI
COWZUQ2hrcK3DvWizvSwC419414gO7WfpZhm1sSatM03RJKzpO5QVAUJmp5z1SeEjk0NL0o3vr3a
dail0qC9ZU+1B5w5mj4R09gwDERKuEa/UohVRXsbmqZUbZ+Cm87fBik/cnqH4I41kpsRME3TC0oq
fdaaYqca9jxDNDUZIR1W4db6jEhUvbAQmGREaj1ua/dVFdmF/oE6n5DMRjSVfc4QjijwJwJJCws1
xMeFlYrEZNtuSG71zF4pnJsgrZ5nK8j8hmlh4ha2EnlD84ibe75rWQEEzGHeai4WorNHIWTkuA62
AbXQPj3gRYeIbeC2JwooMfsU3KpyB3SVdvVq2WyQpbbnvR/oTRfxhSyJLKw067ES/6by29DP2YTz
dS1Sh7JAYIS7TVj4dNci+Ysqvs7g3xKoL3abOHyo+NT+5bYR1LbOIBlIDo1Ai8TacPToLQtksn1/
JQWjelN7eAHS+vlT9b3a3Pi/a61iKD5o9Jp0tSU4wplM7E4ICKwpvYPU20ojeJqbjKb4BMBU9XiR
GwxRN25/LfmulsiUgfBm7nRtGLHhcgPUTBBsibjxoglYAN78we1pPpQunpVxQ55vNK8mP4E5NUGA
G2ZoVWOups4FQ4O8Drxsgnt6natsm+4fxdj9HMMxdhhQA+QOFSJXJh7PgXhZ1R0BZl6zjJaVQ99i
6PR8uVF0behw9nRz5pfj9NMhJdASOy/9hgBmHEQBK4JnpDseGKKq0ZXaf++a7t+Udsh7JNgSWewB
vE6lw95R4ytsU+TbugTQb+kW3r5jpK78ay0HcQapkDUh+A==
`protect end_protected
